//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.02 (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Mon Jul 28 03:25:16 2025

module Gowin_SP (dout, clk, oce, ce, reset, wre, ad, din);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [14:0] ad;
input [15:0] din;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire [26:0] spx9_inst_0_dout_w;
wire [8:0] spx9_inst_0_dout;
wire [26:0] spx9_inst_1_dout_w;
wire [8:0] spx9_inst_1_dout;
wire [26:0] spx9_inst_2_dout_w;
wire [8:0] spx9_inst_2_dout;
wire [26:0] spx9_inst_3_dout_w;
wire [8:0] spx9_inst_3_dout;
wire [26:0] spx9_inst_4_dout_w;
wire [8:0] spx9_inst_4_dout;
wire [26:0] spx9_inst_5_dout_w;
wire [8:0] spx9_inst_5_dout;
wire [26:0] spx9_inst_6_dout_w;
wire [8:0] spx9_inst_6_dout;
wire [26:0] spx9_inst_7_dout_w;
wire [8:0] spx9_inst_7_dout;
wire [30:0] sp_inst_8_dout_w;
wire [9:9] sp_inst_8_dout;
wire [30:0] sp_inst_9_dout_w;
wire [10:10] sp_inst_9_dout;
wire [30:0] sp_inst_10_dout_w;
wire [11:11] sp_inst_10_dout;
wire [30:0] sp_inst_11_dout_w;
wire [12:12] sp_inst_11_dout;
wire [30:0] sp_inst_12_dout_w;
wire [13:13] sp_inst_12_dout;
wire [30:0] sp_inst_13_dout_w;
wire [14:14] sp_inst_13_dout;
wire [30:0] sp_inst_14_dout_w;
wire [15:15] sp_inst_14_dout;
wire [29:0] sp_inst_15_dout_w;
wire [1:0] sp_inst_15_dout;
wire [29:0] sp_inst_16_dout_w;
wire [3:2] sp_inst_16_dout;
wire [29:0] sp_inst_17_dout_w;
wire [5:4] sp_inst_17_dout;
wire [29:0] sp_inst_18_dout_w;
wire [7:6] sp_inst_18_dout;
wire [29:0] sp_inst_19_dout_w;
wire [9:8] sp_inst_19_dout;
wire [29:0] sp_inst_20_dout_w;
wire [11:10] sp_inst_20_dout;
wire [29:0] sp_inst_21_dout_w;
wire [13:12] sp_inst_21_dout;
wire [29:0] sp_inst_22_dout_w;
wire [15:14] sp_inst_22_dout;
wire [23:0] sp_inst_23_dout_w;
wire [7:0] sp_inst_23_dout;
wire [23:0] sp_inst_24_dout_w;
wire [15:8] sp_inst_24_dout;
wire [15:0] sp_inst_25_dout_w;
wire [15:0] sp_inst_25_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_21;
wire mux_o_22;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_45;
wire mux_o_46;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_69;
wire mux_o_70;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_93;
wire mux_o_94;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_117;
wire mux_o_118;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_141;
wire mux_o_142;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_165;
wire mux_o_166;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_189;
wire mux_o_190;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_213;
wire mux_o_214;
wire mux_o_222;
wire mux_o_227;
wire mux_o_235;
wire mux_o_240;
wire mux_o_248;
wire mux_o_253;
wire mux_o_261;
wire mux_o_266;
wire mux_o_274;
wire mux_o_279;
wire mux_o_287;
wire mux_o_292;
wire mux_o_300;
wire mux_o_305;
wire ce_w;
wire gw_vcc;
wire gw_gnd;

assign ce_w = ~wre & ce;
assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_8.INIT = 16'h1000;
LUT5 lut_inst_9 (
  .F(lut_f_9),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_9.INIT = 32'h04000000;
SPX9 spx9_inst_0 (
    .DO({spx9_inst_0_dout_w[26:0],spx9_inst_0_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_0.READ_MODE = 1'b0;
defparam spx9_inst_0.WRITE_MODE = 2'b00;
defparam spx9_inst_0.BIT_WIDTH = 9;
defparam spx9_inst_0.BLK_SEL = 3'b001;
defparam spx9_inst_0.RESET_MODE = "SYNC";
defparam spx9_inst_0.INIT_RAM_00 = 288'h229148A6633198CC6633194CA6532994CA65432190C86432194CA653B1D8EC763B1D8EC7;
defparam spx9_inst_0.INIT_RAM_01 = 288'h33A1D0E87431990C86332190C86432190C86432190C86432190C86432190C8633198CC66;
defparam spx9_inst_0.INIT_RAM_02 = 288'h478BB99ABD5F2F578AC4E271569A4CA65329B4DA7962D371B89C2E07737196B8532150C8;
defparam spx9_inst_0.INIT_RAM_03 = 288'hE4027CFA6C2B08C0C27179A140D78F506C366C36170B84B9DCAE572B1DCADD4C9E4F2772;
defparam spx9_inst_0.INIT_RAM_04 = 288'h3B1DBE6CFD5A9F892271B0942804028584C271F19D38AB4CA2D5EC06DAA534A951A3CFE8;
defparam spx9_inst_0.INIT_RAM_05 = 288'hD2713CA05030184E4735229168B45B329DAF495D9353CAECF2795C6DAE972D98D465B0B7;
defparam spx9_inst_0.INIT_RAM_06 = 288'h32994CA6532994CA6533198CC66432194CA663B1D8EC773B9D8EC7D1F904BE5D26138A06;
defparam spx9_inst_0.INIT_RAM_07 = 288'h432190C86432190C8633198CC86432190C86432190C8643198CC6633198CC6633198CC66;
defparam spx9_inst_0.INIT_RAM_08 = 288'hD4EA71369A4D265329A4D27542D3713C9E4FF7737598C953210EA743A1D4EA743A190C86;
defparam spx9_inst_0.INIT_RAM_09 = 288'h81F9A140D786D06C566C36170B84B9DCAE573BA5CEC15EA6CEE5312703759ABD5F2F97AB;
defparam spx9_inst_0.INIT_RAM_0A = 288'h71B0942804028544C27248F8AA7A4DAAD54AC5E2F176A953240F85D47A00E27F340D44E3;
defparam spx9_inst_0.INIT_RAM_0B = 288'h24124D48A452ADDB2EE794629D72CAEA395CFFCF132786CBE5B0964B0D324EFF621F0943;
defparam spx9_inst_0.INIT_RAM_0C = 288'h229148A6542A194CA663B1D8EE773B9DCEC75389747A3F289BCBA4128944DE5E2E978DE6;
defparam spx9_inst_0.INIT_RAM_0D = 288'h33198CC66432190C86432190C8643218CC6653A190C86331988A45329948A4522914CA65;
defparam spx9_inst_0.INIT_RAM_0E = 288'hB55AB160D271385C2EF77379BCDA5B20CE6743AA150A843A1D0E8753A990C86432190C86;
defparam spx9_inst_0.INIT_RAM_0F = 288'h6C36170B84B9DCAE362B1D8AC15D9DCA22D006FB357ABE5FB3D9CBF572B53A9C4E27158A;
defparam spx9_inst_0.INIT_RAM_10 = 288'h7230DC7C543C26554AA4EAF974984C2953E6350A00E4814615C68181F9A140D786CCAC97;
defparam spx9_inst_0.INIT_RAM_11 = 288'h86CB71E317A75CF4DB9E4F636BA3C15D70F96B853235026A1EC94471B0942804020144C2;
defparam spx9_inst_0.INIT_RAM_12 = 288'h63B1D8EE773B9DCEC7E9BC31646D1E0F49E5F2E9307C5239A00FA5F301C4E4834AA996CC;
defparam spx9_inst_0.INIT_RAM_13 = 288'h432190C8643218CC8653A190C8633198CC66331148A45229148A45229148A6542A194CC6;
defparam spx9_inst_0.INIT_RAM_14 = 288'hF77379BACA5B20CE67442A150A843A1D0E8753A990C6633198CC6633198CC6633198CC66;
defparam spx9_inst_0.INIT_RAM_15 = 288'h0AFD3A99398BC11E4E06FB399CCF6030180C1582BD5EAF5FAC160BE66AF580E1703BDBEE;
defparam spx9_inst_0.INIT_RAM_16 = 288'hC572F954974426552A962A40FE7039230C6181716120D7874CECD86C2E170B84B95CAC36;
defparam spx9_inst_0.INIT_RAM_17 = 288'hDB9EA791B4C8DCAE784B8D7A79126AA30B4571B0942804020102A2723920744B2795D3AC;
defparam spx9_inst_0.INIT_RAM_18 = 288'h6BB5D2DB347CA84B83A1790CE67F2E134BE6E27138A062422554AA66331DB4EF824E6D97;
defparam spx9_inst_0.INIT_RAM_19 = 288'h432190C86432190C86331948A45229148A4532994CA6542A994CC653B1D8EC763B1D8EC7;
defparam spx9_inst_0.INIT_RAM_1A = 288'h442A150A84399CCC87432190C6633198CC6633198CC6633198CC6633198CC66331990C86;
defparam spx9_inst_0.INIT_RAM_1B = 288'h168B45A2D168B4582C258AC562B26134DA4DF6F379BED077375BADE6EB7196B952A110A8;
defparam spx9_inst_0.INIT_RAM_1C = 288'hA5CADD628E3229156581E95900C8874CACB75C2E170B84B95C6C16D9DCA62F057A389C2D;
defparam spx9_inst_0.INIT_RAM_1D = 288'hFA8D46970163234D0481B8D42804020102A261B92492491D904F0AC56AB97AA9431E55ED;
defparam spx9_inst_0.INIT_RAM_1E = 288'h438974984D27980C06F271389C50311CD0694532E192DA763FE2328ADDBF07A6DAE82F54;
defparam spx9_inst_0.INIT_RAM_1F = 288'h331988C45229148A4532994CA6542A194CC6532998EC763B1D8EC76BADDAF189C9DA21CC;
defparam spx9_inst_0.INIT_RAM_20 = 288'h432190EA743A1D0E873399CCC46231188C4633118CC6633198CC6633198CC66332190C86;
defparam spx9_inst_0.INIT_RAM_21 = 288'h469B0986D472B91C6E0773759CDE6E32D96CD6632972A84B219109542A190A843A1D0C87;
defparam spx9_inst_0.INIT_RAM_22 = 288'hA26950FAB67EC86A975C2E170B74B9586C15B94455E6E371B8DC6E371B91C8E47238DA6D;
defparam spx9_inst_0.INIT_RAM_23 = 288'h8238D8280301810282512898745C369749C484CA7960CD531D916AC6738A16DF3FA15449;
defparam spx9_inst_0.INIT_RAM_24 = 288'h02817CBC5E2F940C261422596EC763B1DB0DD78C56735DB8E473B7AA757E72F05C23CD04;
defparam spx9_inst_0.INIT_RAM_25 = 288'h32994CA6532A190C86432994CA753A9D4CA67C2DD2EB77C46632F9C98B90FC4F289BCBA4;
defparam spx9_inst_0.INIT_RAM_26 = 288'h3399CCE46230984C25231188C4522994CA6522914CC66331990C8643198CC46229148A45;
defparam spx9_inst_0.INIT_RAM_27 = 288'h07737598CB652E150BA5CAA152A84B21D12964321D0C863A9D4EA74329D8EC87432150A8;
defparam spx9_inst_0.INIT_RAM_28 = 288'h5BAE170B73B9582BF598ABC9C4E371B91CAF472BD9ECF77B399CCE87BBD9ECF783C1A08F;
defparam spx9_inst_0.INIT_RAM_29 = 288'h512098766F3F9B49832329E93CBE5D259087E6DB0E2D3867A09269F3F184D49475C42876;
defparam spx9_inst_0.INIT_RAM_2A = 288'h0309CD0AA65AAD166B354BBA1B0F8B532FF98ACD2A52F465A44D448238D428030180C282;
defparam spx9_inst_0.INIT_RAM_2B = 288'h432194CA6532994CA61B2E2B55A7CAE170F99D569B132A57938604E2F980DE5E2713C805;
defparam spx9_inst_0.INIT_RAM_2C = 288'h128948A4522914CA6522914CC6633198CC6643A18CC66231148A65329948A6532994CC66;
defparam spx9_inst_0.INIT_RAM_2D = 288'h853A6130984BA213497442612E86431D8EC74329DD10984C25D2C843A1CCE46230980A05;
defparam spx9_inst_0.INIT_RAM_2E = 288'h681381A4E472391CAF5733DDF108843E1F0FB95466351B9549E2B017737198CA5BA952A9;
defparam spx9_inst_0.INIT_RAM_2F = 288'hC20999129C56AE1225D609EDB7538AA8D2483481C0AE8164C3A8565BADD70B74B9582BF5;
defparam spx9_inst_0.INIT_RAM_30 = 288'h663B1588B8684528B49BACDA15097F288FA68238D828030180C2815130A0986E3F1BCA25;
defparam spx9_inst_0.INIT_RAM_31 = 288'h7CAE12E975C365B2D96C2E1B1198C8D09AE8B2697CDE5E2F13C805130184E68552AD1449;
defparam spx9_inst_0.INIT_RAM_32 = 288'h128944A4522994CA65231188C4623118CC6623AA18EA642A190E685421C8E2632A954A85;
defparam spx9_inst_0.INIT_RAM_33 = 288'h94CA612E8744A210E863BA2110984C25D2C864A24D0472391C4FE6130944A25229148A45;
defparam spx9_inst_0.INIT_RAM_34 = 288'h884C6A572B95CB27D4EA7536973B9E4E64B03783B99ACA53A550A8854AA554AA552A954A;
defparam spx9_inst_0.INIT_RAM_35 = 288'h343A79929A98BFCE2965E988CA6F5542A2352B1DD2EB73B8572731682BD1E8E4723D9EF0;
defparam spx9_inst_0.INIT_RAM_36 = 288'h2914821CE17A4315C3A2C91C6A24120902616138A87A51311C0DC5E2F17CA88A562A90E6;
defparam spx9_inst_0.INIT_RAM_37 = 288'h6C365F2F97CBE5B2D888E2C4BE51309BCBC5E27100C6844A2110A9253B1D86A354BB1F4E;
defparam spx9_inst_0.INIT_RAM_38 = 288'h231188C4623198CC6633998CC654329D90E9743A59087432150A644BAE1B0D86C2E170B8;
defparam spx9_inst_0.INIT_RAM_39 = 288'h74422532984C25D2E964AA4D0482391C4E27230984A25229148A45128944A45229148A45;
defparam spx9_inst_0.INIT_RAM_3A = 288'h0AFD7A993C9ED2E711378BB998CA53A590E9854AA976BB5DAED54AB562A95088442210E8;
defparam spx9_inst_0.INIT_RAM_3B = 288'h559A40C86B49B724152B1592E973B057677288BC15E8F4723D9EF0784C6A592D9F53E815;
defparam spx9_inst_0.INIT_RAM_3C = 288'hC2D1206C26128542816138A47A51311C8C06E2F174BC433D2692C654B25516BF6C4F1AAA;
defparam spx9_inst_0.INIT_RAM_3D = 288'h8C9DA638B02D0B062602F13CA4754A2490471492494492522D58CCA75BA9B0BB67B69466;
defparam spx9_inst_0.INIT_RAM_3E = 288'h641988A8673BA2136BD5FB3DB8B9439D4C655BAE1B0D85C2E130B86C361B0D86C361B2D9;
defparam spx9_inst_0.INIT_RAM_3F = 288'h54AA510682391CCE68339184C26231188A45020104A25129148A45231188C4633198CC66;

SPX9 spx9_inst_1 (
    .DO({spx9_inst_1_dout_w[26:0],spx9_inst_1_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_1.READ_MODE = 1'b0;
defparam spx9_inst_1.WRITE_MODE = 2'b00;
defparam spx9_inst_1.BIT_WIDTH = 9;
defparam spx9_inst_1.BLK_SEL = 3'b001;
defparam spx9_inst_1.RESET_MODE = "SYNC";
defparam spx9_inst_1.INIT_RAM_00 = 288'h4813BDB8BA54261329854AAD78CD66B3176BB562ED52984CA6530874426532984B2190C8;
defparam spx9_inst_1.INIT_RAM_01 = 288'h1B158EE973B0D7E9B3B94C5E0AF47ABD9EF0784C725D3FA0546A560AFD76973B9E52E732;
defparam spx9_inst_1.INIT_RAM_02 = 288'h6138A47A41319CCE47F289B8B43F2CA755284411C8DACB5C49622824B2C0CA8A4F2F67D4;
defparam spx9_inst_1.INIT_RAM_03 = 288'h02F978BC5D2F99132B2481FCE2914FA3D24A35AAD96EB95D2E14C9E2E12870270B8582C1;
defparam spx9_inst_1.INIT_RAM_04 = 288'h57D4726F106E2A12A75BAE170B84BA5D2E986C2E170B85C361B0F96C4663297B98B54F83;
defparam spx9_inst_1.INIT_RAM_05 = 288'h4419C8E4623198CC46120904824120904824231188C4623118CC66531150D29B552AD7ED;
defparam spx9_inst_1.INIT_RAM_06 = 288'h9552F19CDF6FB399ABB56AF99CBE5F33598B84C2653296421D0EA7542A150872391D10A8;
defparam spx9_inst_1.INIT_RAM_07 = 288'hEA64EA4F067ABDA0F09854765F40A0D46A35EAED32973A9CCA24D15813FDB8BA54261329;
defparam spx9_inst_1.INIT_RAM_08 = 288'h1291BCB43C221E958A541199129C5EB2A92BF422890C9A50B725B31B158EE973B9586A15;
defparam spx9_inst_1.INIT_RAM_09 = 288'h752205008F469F9029048A9570C963A952A902F13074290C0602E18140A87A41299CCE67;
defparam spx9_inst_1.INIT_RAM_0A = 288'h3BA5D2E974BA5D2EB85C2E130974C2E1B0F95C2DD2EB78CBE3662C128140BE6F30189089;
defparam spx9_inst_1.INIT_RAM_0B = 288'h128904804020104824229148A45229148C460211613CDE6DAED7ED98FD06D944873254A9;
defparam spx9_inst_1.INIT_RAM_0C = 288'hE59355EAF57ABD1E4EB54A613096421CCEA743A2150883399D50C964AA10E6733998CC66;
defparam spx9_inst_1.INIT_RAM_0D = 288'h9854725D30A0D46A15DA6532773993451E4F270BBDB8BA5526D56AB5E3399ED06837D9CC;
defparam spx9_inst_1.INIT_RAM_0E = 288'h84CA9D2A794B2265B555925546995AC223D31B1592EB74BA5CEC761AFD32751883C1E110;
defparam spx9_inst_1.INIT_RAM_0F = 288'hF47A0528A559A4504812F934762B0D064321A1D0EC7C412998CC66128178B6491D0C0CE8;
defparam spx9_inst_1.INIT_RAM_10 = 288'h5C2E12E974BAE170D85C36170763B3DE30D7988B54FC4E20184C0684C2913E7C369F91E8;
defparam spx9_inst_1.INIT_RAM_11 = 288'h128944A25129148A45434279A50F7C2D52C94754B26B1E6D2DD2682B158EE974BA5D70D8;
defparam spx9_inst_1.INIT_RAM_12 = 288'hF6DA9D2E974AA10EC843A1D50A8542A190E974B2590A853A9D0C66229144804020104824;
defparam spx9_inst_1.INIT_RAM_13 = 288'hDA64F27738923C5DEDE67B7DBCCD5EAF97CBE6733D9ECF67B3D9EC162BE211178B41604F;
defparam spx9_inst_1.INIT_RAM_14 = 288'h082AD9628751C15FF40A9592EB85BA5D2E972B0D7A992A8CC62311984C2E3B2FA0502A14;
defparam spx9_inst_1.INIT_RAM_15 = 288'h1301789A3C160AC562C1E0F47E4232190C6643097CBA591A8605C543EB2138B74322D794;
defparam spx9_inst_1.INIT_RAM_16 = 288'h3BB6675195BA592C96ACADEA38A12F13CA2653BA59207B2E1B4FA6F47234FE8048A4928A;
defparam spx9_inst_1.INIT_RAM_17 = 288'h95734A072F84B0D027B47B3D909231184DE60A8D8EE975C2E170D85C2E170974BA6170B8;
defparam spx9_inst_1.INIT_RAM_18 = 288'h43A9D50C884C26130985425D2E97431D0E66329144804020104824020104825128944A25;
defparam spx9_inst_1.INIT_RAM_19 = 288'hC67B45C0DF67B019EB06FB399CBE5F2F97EC06239E0F058240DE2F275AD90C874B2150C8;
defparam spx9_inst_1.INIT_RAM_1A = 288'hFA8D92EB85BA5D2E973B0D429D3C954AA331A8542A392E9FD3E9F4DA5CEA5527813BDBEC;
defparam spx9_inst_1.INIT_RAM_1B = 288'hE2713C8455331D4E864311BCBA5A238DC503C1A9E95ECB562D51CC695B5146A75EB55FD3;
defparam spx9_inst_1.INIT_RAM_1C = 288'h0A35EB2B6A87290DC302219D2C903D96CBA6E47A391A7E40A516AB2401FCBC4D1E8F47A3;
defparam spx9_inst_1.INIT_RAM_1D = 288'h3239D4DA39058B87A40A8D92EB86C2E170B86C2E170B85C2E130989D360EE764B258EC76;
defparam spx9_inst_1.INIT_RAM_1E = 288'h95426130984B214E66329144A24020104824020100804020940A05956B4625208EBE98C9;
defparam spx9_inst_1.INIT_RAM_1F = 288'h1683397ABC56AB97EB16239A0B0479BCDE4F37DAD0EA8643214EC85429D90E99552A5509;
defparam spx9_inst_1.INIT_RAM_20 = 288'h3B1582BF4D9DCAA551C8DC6E392D974FA7B3C9D4A63115783799ECE60B8DE4E06833D7CB;
defparam spx9_inst_1.INIT_RAM_21 = 288'h228978B44A2E1648A190D06D529068BB994A5973C52EC96C2DA192EA0D92EB85BA5CEC97;
defparam spx9_inst_1.INIT_RAM_22 = 288'hE109213AC75E1A8BC7B372011C7E3824D46A248A3CDE5F279389C4E27900A6663BA1CEC7;
defparam spx9_inst_1.INIT_RAM_23 = 288'h0A9592ED86C2E170B86C361B0D85C2E12E975C1DCEED86C1D86A555B15426345A9511AE7;
defparam spx9_inst_1.INIT_RAM_24 = 288'h12998CA04F180C060332687022463DAAD6EB95E36DB6EF80439FAFA59A3CBA4D1D86C3A2;
defparam spx9_inst_1.INIT_RAM_25 = 288'hE59B59C8E268B49C4F16DA950A864A2150E995426536AD5EAF174A94CA612E87431D0C65;
defparam spx9_inst_1.INIT_RAM_26 = 288'hC964B2592D96CFA7D3C9545DE8D16030182D27138DC4D16830180C1603397AAC4EA755CA;
defparam spx9_inst_1.INIT_RAM_27 = 288'h61A0AC94A26F2F564DC5D2DD6CC65AAB9BD4C91D9AE763B35DAE963B1586A14EA6CF2572;
defparam spx9_inst_1.INIT_RAM_28 = 288'hE2E9B4FC8D469FCE48B38A491E6028940A05129150CC7843A18EA732897C984B1C8DC6A2;
defparam spx9_inst_1.INIT_RAM_29 = 288'h4BADD6ED86C2DD2E973B9D8EC963A9D4A85409FCBE5F219954EC963621784C7A519EC964;
defparam spx9_inst_1.INIT_RAM_2A = 288'hE1915D18B26A3C9FEE2793F1AAA5532E59AED6BA80DA4A140685C43B2592EB75BAE16EB7;
defparam spx9_inst_1.INIT_RAM_2B = 288'hF652950C964B25D32AB5D2A556AC5EAF176AA54A610E863B1D0C65230940804120904804;
defparam spx9_inst_1.INIT_RAM_2C = 288'h983BD1A4C160B0580C168B45A2D168B0180C05FAF95CAD56A753CAD50B11A6D260B45C2E;
defparam spx9_inst_1.INIT_RAM_2D = 288'hC5DADD6AB451A6D932FA0D4EC964B2DD6E963B1D8AA14FA74F65B2D96CB2592C964B65B2;
defparam spx9_inst_1.INIT_RAM_2E = 288'h148238C0734017886632A194CE794421D0C743117C9A4B1C8DC6C251A060446B57B399AB;
defparam spx9_inst_1.INIT_RAM_2F = 288'h2B158AC552A0CC2412D96C7A5D2099512AB67BECA9181125AA136481E9BCF87D412493C6;
defparam spx9_inst_1.INIT_RAM_30 = 288'hD9F5625CE658238E08F3F984E671369287842B1D92EB75BADD2E974BA5D6EB75BA58EC76;
defparam spx9_inst_1.INIT_RAM_31 = 288'hE66AED78BC5EAF578BA54A610C763A990C854301386242281387E4F2D2C1C4F681BFDC50;
defparam spx9_inst_1.INIT_RAM_32 = 288'h371385A2D26934580BF57ABD5CAE56A753A9B4F28564C260B019ECB5C2590E974BA655AB;
defparam spx9_inst_1.INIT_RAM_33 = 288'h0A74C28965B9D8EC963B1D8AA350A7D3A7D3FA74FA7B2C95C6E3718833D1A8D5733D5C6E;
defparam spx9_inst_1.INIT_RAM_34 = 288'h6331DCF28A4D2610E853197C9A3B1C8E06E2613094322336AFD94AA552DD4AA45121D22E;
defparam spx9_inst_1.INIT_RAM_35 = 288'hD8EC7A3D1E97CCA8954B3DCE8AD52F8D0F6AD3391C7C7349A4926975A2811E7349204C87;
defparam spx9_inst_1.INIT_RAM_36 = 288'h71D10D1CD17736990C2B1D92CB75BADD2E975BA5D2E963B158AA552A954A83409FCBA3D1;
defparam spx9_inst_1.INIT_RAM_37 = 288'hB54A5D0A7532190C8532F8C066522E8F8666F73C9A49138632D7121AA5BAA90A679E06C2;
defparam spx9_inst_1.INIT_RAM_38 = 288'hF57ABD5C9E4EA71388C46A7D40A05FAF556974321910984C26D5CBF6F3399CCE6733176A;
defparam spx9_inst_1.INIT_RAM_39 = 288'h2A954AA351A0D46A351A8D429D3D9646A150B8D426150B8E4AE57188B411E8E47234980B;
defparam spx9_inst_1.INIT_RAM_3A = 288'h63A1809A3B1D0E470281C0942A0D1C27DBEDA552DD4CA75A24D0EAA96CC28764B1D4EA76;
defparam spx9_inst_1.INIT_RAM_3B = 288'h2B0D16B37D8C9C48A6555958585138A0D30C8673E5BE804329D2A8944A29169B4DA65308;
defparam spx9_inst_1.INIT_RAM_3C = 288'h2A958EC965BADDB0D86BADD2E762A9546A343A95027D2D8EC763D1E97C825D1D8EC7E434;
defparam spx9_inst_1.INIT_RAM_3D = 288'h2209088850268D4E4EBA550E210D691C8EB0D95C85AA8E3511C7248240F08C9E693CE2B2;
defparam spx9_inst_1.INIT_RAM_3E = 288'hC462311A9D4DA20CE663B1DD108944A2D3CBF67B01A0D06733176AA4CA18EA6432150A85;
defparam spx9_inst_1.INIT_RAM_3F = 288'h4B1D8AA34F9ECB2350C96CBE7F3E9F4FE814EA64E62F067AB8DA2C258AC15CAD4EA71188;

SPX9 spx9_inst_2 (
    .DO({spx9_inst_2_dout_w[26:0],spx9_inst_2_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_2.READ_MODE = 1'b0;
defparam spx9_inst_2.WRITE_MODE = 2'b00;
defparam spx9_inst_2.BIT_WIDTH = 9;
defparam spx9_inst_2.BLK_SEL = 3'b001;
defparam spx9_inst_2.RESET_MODE = "SYNC";
defparam spx9_inst_2.INIT_RAM_00 = 288'hA1C89C4E191016D68F16FB696EA85B28906816D48AA552A9D4EC552A15068342A9D4EC96;
defparam spx9_inst_2.INIT_RAM_01 = 288'h24328D12260F99D70CB69C862AB24A29950AB4DA6D38AC55A6932863A184BC4C1D8E8543;
defparam spx9_inst_2.INIT_RAM_02 = 288'h6BADD2C752A8D068131984B6370B864363F1098CC67F2D8E47A5F33B15468544A7479403;
defparam spx9_inst_2.INIT_RAM_03 = 288'hEA3CC21CFB6F1B08EA36EAC4AA13020545035118183E474DAF1BAE2A954AA764B2DDF0F8;
defparam spx9_inst_2.INIT_RAM_04 = 288'h8349E9168B4522D389E5F33D80CF672ED5499439D8C8642A150A8542990CA6501893D9F4;
defparam spx9_inst_2.INIT_RAM_05 = 288'hC974C2814FA75028351B7D6E7318833D1C4D469B4980BF572793C9D4E22D168A3C19CAE4;
defparam spx9_inst_2.INIT_RAM_06 = 288'h782BF992A95BAD126994B402834F9954EC352A0D068342A9D96CD75BADD2C751A7CFA5B1;
defparam spx9_inst_2.INIT_RAM_07 = 288'h28A492451C71A4914BC562B158AC55A6912863A184BE4E1E8F0762B1C8A854380D090E2D;
defparam spx9_inst_2.INIT_RAM_08 = 288'hD863EDF4EA7E43A213098D0683309FCFE614E99D4EA141A1D7A4AD02B21D3E570C8D5410;
defparam spx9_inst_2.INIT_RAM_09 = 288'h4311A866020184828120B88CE2D8823F1AEB1A8D4AA563B25D6ED74B254EA5409FCFE5D2;
defparam spx9_inst_2.INIT_RAM_0A = 288'hC56AF97CBD5E2A932883B1D4C8542A954A8552A14CA641219755306883F5FF1F8CB49207;
defparam spx9_inst_2.INIT_RAM_0B = 288'hFAED2E7327833D5CAE572B91C6D260AC140AF4EA6D168A3C9A8D87D3F1F91C9D4EA71369;
defparam spx9_inst_2.INIT_RAM_0C = 288'h547B2A3D3F98506A553A150A8542A9D92CB75BADD6E963A8D027F3C96CFE9F4FA7D02A35;
defparam spx9_inst_2.INIT_RAM_0D = 288'hC5E2AD58AC4DA24F0753A188A04F270F4782B1D8F07A4B1487C8E716A3C5D8CB5C2D548A;
defparam spx9_inst_2.INIT_RAM_0E = 288'h0A0D0AA553A9546A352A04FA8355BADCE8333641CCCA8F330B4DCE7A45269B68A53490CA;
defparam spx9_inst_2.INIT_RAM_0F = 288'h106141A769C0549F2CFA050AA763B1D8AA351A0D02613E96C7217096D369D6FD8FC82634;
defparam spx9_inst_2.INIT_RAM_10 = 288'h73B194C8552A954A8542A10C885321114D281379854EED87C5DB8680489424040A8904C2;
defparam spx9_inst_2.INIT_RAM_11 = 288'h57ABD9ECE57230962B157A753A9D4E239049138A092290572B1368B4E2B158AB4DA69128;
defparam spx9_inst_2.INIT_RAM_12 = 288'h4A9D0A8542A9D52C965B2DD6CB64B1546814D9ECFA9D4FA8D46A35CA5D2A711682BD5ECF;
defparam spx9_inst_2.INIT_RAM_13 = 288'h532188A240278F87A3C1E8F89C4D1E0B05A253FB0DC0DD6CAD548A43D291D92F9F4C2876;
defparam spx9_inst_2.INIT_RAM_14 = 288'h5A3DDB036EAFD0A894AB2B50C4613D120786AAEDC2E380BA459608C5E2AD569B4D224F06;
defparam spx9_inst_2.INIT_RAM_15 = 288'hD9FD0AA964B0D7E9B3E974BA5D1D85BE9F2E864B6DDD009150EA751A954AA964B258AA35;
defparam spx9_inst_2.INIT_RAM_16 = 288'h32B198C8532A18CA04A1D12CBC8F4F230F8671F99502580980C2A4106909A53D8F2A540F;
defparam spx9_inst_2.INIT_RAM_17 = 288'h2602FD5E9E3E9B8C070309C5009F4EA351A8C4E271389B4D225107833998CA552A954AA5;
defparam spx9_inst_2.INIT_RAM_18 = 288'h3BA5D30B85C25CAC15FAF576BD5FB7DBAB9479345A0F078341A0F098CC6611077B395C8D;
defparam spx9_inst_2.INIT_RAM_19 = 288'hE2F1349A4D1F13C9E422F2D1C0DD67BADA6A251265551B8A556EB76C361B0B74B9D8EC76;
defparam spx9_inst_2.INIT_RAM_1A = 288'hF92D2DF6773A1ECAA39224974791C6581ECA65E371749D4DA1CCC6532148A451281009E4;
defparam spx9_inst_2.INIT_RAM_1B = 288'hE96C763B0A7431D90CA75BF62121A154EA754B2592C963B1D4EA755BADD6C962A8D02814;
defparam spx9_inst_2.INIT_RAM_1C = 288'hA1C09C70592C114682A22209D3278FB9D66A50C8DD26DE50138AEB098502613F9F4BA5B2;
defparam spx9_inst_2.INIT_RAM_1D = 288'h13920924A1502BD5EAE5F2F97CBD562AD349A45224F0773399CCE642A990A6542A148A04;
defparam spx9_inst_2.INIT_RAM_1E = 288'h0B7D7AB94AA4CE2512489C09E6F47ABDE151C9E4F6792A8C3D5C8D4692C1409E469F8E08;
defparam spx9_inst_2.INIT_RAM_1F = 288'hE1B1FD66E3703A988A250A2144DC8955F0F97CC6632F85C25CEC563B9DD2E975C2DD2E76;
defparam spx9_inst_2.INIT_RAM_20 = 288'h81F1DA6DBFC5D669AE44A27160CA439A0F06532148A251281009E4F2F1749A4D2713C804;
defparam spx9_inst_2.INIT_RAM_21 = 288'hB8647E4332A9D52C964B2592C964B2592CB64B2DD6E963A9546A345B647E5B1A4094CFC6;
defparam spx9_inst_2.INIT_RAM_22 = 288'h40693DA369D1E2687175920D0C802382C8ECF9FCFE7D2E96CB63B1D8DC2DF4E86BB2194D;
defparam spx9_inst_2.INIT_RAM_23 = 288'h168B45A2D06833D9CCF5F2F5589B4CA2512873A990AA653214CA6502D8D84A261A888020;
defparam spx9_inst_2.INIT_RAM_24 = 288'hF76B719CC069B9E172D9F4FA9D3C94415C6D569B0962A04FA0104945AAD9AAD469B49A4C;
defparam spx9_inst_2.INIT_RAM_25 = 288'h35021534AE9955F0D87CC6675396C25CAC354B9DCEE974BADD6E972B0DBAB53488BC1E0F;
defparam spx9_inst_2.INIT_RAM_26 = 288'h9601E562D8431AD0E653218CA451289009E4F2F9389A4D1F0FC803E2012104D678B6D92C;
defparam spx9_inst_2.INIT_RAM_27 = 288'h4B258EC552A9D4EC964B25D6EB74B1D8AA553A9506833A85248CC8B2984D5B71CFDEEA50;
defparam spx9_inst_2.INIT_RAM_28 = 288'h598C79D4B44018910DF9FCFA7D2E974B63B1B7CB9DAEC763B29DB0D974BE6343AA596CB7;
defparam spx9_inst_2.INIT_RAM_29 = 288'h371B89A0DF672F578AC54A1CF0773A998D088401604C2613090060101038A0EBA5D1A691;
defparam spx9_inst_2.INIT_RAM_2A = 288'hD9ED3A9B3C94C59EAE66A34D84B158A894AC874BE61308834160B057ABD5EAF47A3CDE6E;
defparam spx9_inst_2.INIT_RAM_2B = 288'h6C3E675397C25C6A154B9DCAC563B25D2E973B8DB6AF217E36592B652A55129C58B59F51;
defparam spx9_inst_2.INIT_RAM_2C = 288'h63298CA452289409E40279389A3D1F0FC60323010CB8A2683399ED659A44EC9DA25D7097;
defparam spx9_inst_2.INIT_RAM_2D = 288'h4B2DDAED75BA58EC75FA35CABD23A5C690861459606EBFBA6A685038B29534A844A2D0C5;
defparam spx9_inst_2.INIT_RAM_2E = 288'hFA7D3E9F3F9F47619096BB196CC764BB21F2D9F5028353B1D92C966BAD8EA551A8D4AA76;
defparam spx9_inst_2.INIT_RAM_2F = 288'h0672F15698431A11AAC599E46A1512850060401018206753A994EBC71456651E74B09346;
defparam spx9_inst_2.INIT_RAM_30 = 288'h672B91A8D3612CD6CC87CC2A352A94CA65328944A251288BC5E2F178B41A0AF371385A0D;
defparam spx9_inst_2.INIT_RAM_31 = 288'h2B0D42A351B158AE570B6D66691F75315248F2F944CE8C58B5A152EA7D3A9D3C954620EF;
defparam spx9_inst_2.INIT_RAM_32 = 288'hF278F87C3E1F8C060353994CAE7B4F2F99CDA642F8C8858AE130D86CC6675396C1D82BF4;
defparam spx9_inst_2.INIT_RAM_33 = 288'h1AF50AA35E91D76307441A20704D7863AC9128E39122784E2A8F0673B190A65329144804;
defparam spx9_inst_2.INIT_RAM_34 = 288'h863AD970DA75C36213FA7D46A553B1D8EC755AA54EA541A154EA764BADDB0D75B9D8EA55;
defparam spx9_inst_2.INIT_RAM_35 = 288'hC599E88C361A88C04051285C564D2D928965D3AAE9D0C551A68A00E9FD02813F9EC6DF2E;
defparam spx9_inst_2.INIT_RAM_36 = 288'h5733E2352B9DCEE994BA5D2E753A9D4E6733994CA251178B41608F371345BEBB4CA293AB;
defparam spx9_inst_2.INIT_RAM_37 = 288'hBA448E1EEB63A88FC5B1E0C4B08F61BA2172EA6D36793B94C620EF77B3D9EAE469B0D8AC;
defparam spx9_inst_2.INIT_RAM_38 = 288'h4329D8CC69462B174AD6DB38C2795FD9313A8D4EA75196C15829F3FA7D02A151B05BEBD5;
defparam spx9_inst_2.INIT_RAM_39 = 288'h8411BCD03820C0F354B6EB9940764D264F8883B9D8C85429948A2401F8FC7E3F180C4844;
defparam spx9_inst_2.INIT_RAM_3A = 288'h1A8D4EC964B1D4EA55F97CBE5F2098D0AA754BADD6EB74B1D8AA551A0502A150A0D46991;
defparam spx9_inst_2.INIT_RAM_3B = 288'h0090542E170B89C6E4825168B058238D4420C96CFA7F3E95C25CED863AE194EC86C7A614;
defparam spx9_inst_2.INIT_RAM_3C = 288'hEAED76994BA5CEE773A9D4EA753A9CCA2512683415E4D0672F15495479A8B2592B914460;
defparam spx9_inst_2.INIT_RAM_3D = 288'hD1F8CCB49F61B9A131A95CAE572A8CC1DEEF572395ECF572351ACD5733E2152B9E4F29B4;
defparam spx9_inst_2.INIT_RAM_3E = 288'hD663194271413C6CF87CBE5F2D84B15468141A8D4AC560B6D264D1380BF9D4B5489B8983;
defparam spx9_inst_2.INIT_RAM_3F = 288'h28639968934322916893C1DCCA653214CA451188C0604121110A854331E5148A4526954A;

SPX9 spx9_inst_3 (
    .DO({spx9_inst_3_dout_w[26:0],spx9_inst_3_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_3.READ_MODE = 1'b0;
defparam spx9_inst_3.WRITE_MODE = 2'b00;
defparam spx9_inst_3.BIT_WIDTH = 9;
defparam spx9_inst_3.BLK_SEL = 3'b001;
defparam spx9_inst_3.RESET_MODE = "SYNC";
defparam spx9_inst_3.INIT_RAM_00 = 288'hC7EC361D1F90CCA8743B2592C963B1D4AA75F9AD86BF45B8D766F777C20CFC64179D65D6;
defparam spx9_inst_3.INIT_RAM_01 = 288'h91A88C4A361A0502C3C964B65B2C8DC25F0EA6CB25B8FE8F4BE7F41A9552C964A9D06613;
defparam spx9_inst_3.INIT_RAM_02 = 288'hA9D4EE774B9DCEA7539954A22AF57A3B98E8D2D120926B3C95868100884802020285C6E4;
defparam spx9_inst_3.INIT_RAM_03 = 288'h88CC6E5B3D964AA330269391CCF67B39DD0E77C42A392C9E4F2994FB7576B95CA5D2E974;
defparam spx9_inst_3.INIT_RAM_04 = 288'h4BA5D2E762B154A8554B2DD6E970AD4D21EEE76B698A903612C762020914D49E58B0DCAF;
defparam spx9_inst_3.INIT_RAM_05 = 288'hA449DCEC653218CA45220904824221954AC673C1ED3AAC4C2255ACB5DAFDC48F3BAB6835;
defparam spx9_inst_3.INIT_RAM_06 = 288'h2A9D4EC753A9D4EA952A0D16CB80B158EFB38B2B90E27D320BCF951BE3554CA13A1F1306;
defparam spx9_inst_3.INIT_RAM_07 = 288'hC964B2391B8DC2DF6FB6CB69D90E8FCBA7F41A154EA953A8D3E5B1E87C02212299D0E894;
defparam spx9_inst_3.INIT_RAM_08 = 288'hBAD566913893C49DAC03B8E07249251144410010482201018584E36138D848140A8584A1;
defparam spx9_inst_3.INIT_RAM_09 = 288'hD74B061769A2C9A49157ABA6170985C76572D9E4EE75399D4EA75398D4B2793B9D4EE994;
defparam spx9_inst_3.INIT_RAM_0A = 288'h4C260F037DABC81D8CC64291006D260F07C343117158AC57B3DB52FB9E5F73C6D85E2651;
defparam spx9_inst_3.INIT_RAM_0B = 288'h321950A85532998EC794DA713AAD562B158B655AFD98B3401E96F0D8EC7A4141A8D4ECB7;
defparam spx9_inst_3.INIT_RAM_0C = 288'h2A154AA763B154AA550A35EA0E6026964B88FC3D1572C3481BDA67C3D9E8EE6429954AE5;
defparam spx9_inst_3.INIT_RAM_0D = 288'hD8642E191D97CC2613FA8D8EA74197C7E211299D12A953A9D96CD73B0D46A562B0D4AA76;
defparam spx9_inst_3.INIT_RAM_0E = 288'h2438DC6E361C0D024110884000000209C7035130984A240A894261C85C2E151B8DC6E16F;
defparam spx9_inst_3.INIT_RAM_0F = 288'h268B51ACE56BBA613098CC663329954EA753A95CEE7529944A6754BADD6A953A9CC9602E;
defparam spx9_inst_3.INIT_RAM_10 = 288'h752204DE5E268FC82542C1F1549F664CEEF9BEEFB7CDAAA7399669E3719D7F028AC965EF;
defparam spx9_inst_3.INIT_RAM_11 = 288'hB562B95CAE56AB158A84DAB574A3401D53AC8743AA191D974C6A976CAE0F057FB4CC5D4B;
defparam spx9_inst_3.INIT_RAM_12 = 288'h6C0D426CE32E138F26A6D54626A34AA9D4C9D459E8D06733198CC542A154AC673C225149;
defparam spx9_inst_3.INIT_RAM_13 = 288'hFA0502611E8743E0114A2556CB64B2596CD73A954AA752A8D028341A0D0AA553B1D92C96;
defparam spx9_inst_3.INIT_RAM_14 = 288'h21084000020C0ECB6561B0D4461209850261A753EA171C964763B0C86432190E8FC82412;
defparam spx9_inst_3.INIT_RAM_15 = 288'h5733DE132B9E5329B5B9DCEA51168341E533BADD6EB74BA5D2249065491C6A25130CC261;
defparam spx9_inst_3.INIT_RAM_16 = 288'h83EAB15ECB9CEFFFFFFFD77AC92181C5E7349A1435D2C65DB46271F6FB0D88C259B1DCEF;
defparam spx9_inst_3.INIT_RAM_17 = 288'hB45AAD72B5491C9089462B61F70C8EC86AB76CA60EE570B54C1D2B5419C0A0402090CAC6;
defparam spx9_inst_3.INIT_RAM_18 = 288'h92042690C353284EC9C4DA2CF46A3C9E0CC5633198CE783CA2D38AC56AB95EAE4F2753A9;
defparam spx9_inst_3.INIT_RAM_19 = 288'h5AB59EED76BADD6EB74B154AA551A7CB65D20984C68553B2596EB76CFD4EA34F58978B45;
defparam spx9_inst_3.INIT_RAM_1A = 288'hC3595C66120A0944A286CBEA192E974BE5D1C864321B0E884423F1097C7E1CFD773C6273;
defparam spx9_inst_3.INIT_RAM_1B = 288'hEAE52A4F04723DA112AA552E974CA5D226B195D11C6C25138D04A231188824151D178DE7;
defparam spx9_inst_3.INIT_RAM_1C = 288'hEB5D6ABD64D5733D9EEF47174388A6BE1AEDA5DA856AC25128D86C26235DF52DA7D42C16;
defparam spx9_inst_3.INIT_RAM_1D = 288'h059B21D90D86C82AB86CAE170981B54C9D6B94B210C8642A95CD48E57AF15B3BDF7BFFBE;
defparam spx9_inst_3.INIT_RAM_1E = 288'h84D230FA7C3D1E4CE683C19CCE783CA2D38AB562B95CAE4F2793C9D3E26D76C95B24D029;
defparam spx9_inst_3.INIT_RAM_1F = 288'h4A9502612E8E42DF90F97C866543AA592C960B1DC6A34E9EAB49E5B269820B3868A45068;
defparam spx9_inst_3.INIT_RAM_20 = 288'h86D3F23F30A0502612D8EC761AFE7FBF9FCFE7F3F5DADD77BCA4936B359EEF77BB5D6EB6;
defparam spx9_inst_3.INIT_RAM_21 = 288'hAA5D32994CADD666B2A651184C26138D44C241B0DC8C3725170DA6F3F1F0D0471B8DC6E3;
defparam spx9_inst_3.INIT_RAM_22 = 288'h8E677BDFECEFE31FC9E311B126B350A415CA151B1DF72EA858AE57FB756A4CF369B55F11;
defparam spx9_inst_3.INIT_RAM_23 = 288'h4BAE1B0B82B5CD1E0DC5D26110783C1A91A9159311F3AFFFFE7BF8697DEBBFFFFEFB3B9E;
defparam spx9_inst_3.INIT_RAM_24 = 288'h93C1E0F079452715AAC56AB55A9D4E2311A8D36A7578CC5CA9542994F295B6FC7DC36615;
defparam spx9_inst_3.INIT_RAM_25 = 288'hE8FC868754AA58EA55FA9D828134ACC21065F330BCE93189A892084442311C8D3D1E4D27;
defparam spx9_inst_3.INIT_RAM_26 = 288'hE9747A1CFE7F3F5F8FC763B5DAEE7840A4946B3DDEF188C35D6C9619FCB6390B7D3ADF8F;
defparam spx9_inst_3.INIT_RAM_27 = 288'hA651144A25130D02A251C124B0471B8E0703A2E1B0D459238D4461A7E43E6352A8D46833;
defparam spx9_inst_3.INIT_RAM_28 = 288'h51C8D8C49551A455C90492D9D51EA0586E570BF56A2AE261315F11B9E536BB5DAED6A8F3;
defparam spx9_inst_3.INIT_RAM_29 = 288'hF5EA6D168B4623520AE53382BDDFFE78B2F47DD777DBEBED773DDF9E77AF8DADEDF969A9;
defparam spx9_inst_3.INIT_RAM_2A = 288'hF5FAFD7CAC4DA2CF67E472795ABC5DAD9449344A4972DB753EE393FA0D4EC55FA5455C6D;
defparam spx9_inst_3.INIT_RAM_2B = 288'h3B74C6875F97CA1F0702F95C68B49E3CD42803AA313C9D451E8F6783C1E4F48B4EAB960C;
defparam spx9_inst_3.INIT_RAM_2C = 288'h088446231291CD28B56BB5DEEF77BB592A74D85BE5D4EA753B1FD0E8FC866543A1506833;
defparam spx9_inst_3.INIT_RAM_2D = 288'h51B91C8E361B8D84A25138DC6C361288C220C8FC8AA763B154683409FCBE1CFF7FC3E3D2;
defparam spx9_inst_3.INIT_RAM_2E = 288'h141A99D51DA0542C370C6D6628D159315F11B9ED3ABD5EB6DAEB34D759544A251288C2A2;
defparam spx9_inst_3.INIT_RAM_2F = 288'h05B3D71DECF16AADB7BED76BB9EFFFFFBF7DBEFFB395BEF2EEDEE621A848A29652A8D40A;
defparam spx9_inst_3.INIT_RAM_30 = 288'hE57275188D56AE1468042A794CCA6D3AA172C964B65B2C8CBD9C8D15FAB93C9E4F28166C;
defparam spx9_inst_3.INIT_RAM_31 = 288'h642230B25969499669E39A293AAD4E22CF6793C9E9169C572FD80C0582FD7EAE56A753A9;
defparam spx9_inst_3.INIT_RAM_32 = 288'h4B2592CB65A9D025B1C7D3A5B4EB7536DDAFD86C3A3D1F97CBE5F22A7446653C8747A4AD;
defparam spx9_inst_3.INIT_RAM_33 = 288'h6130D446130A0544A2D9050EC973B9586A54F97C7A1F00894CEA765B2D96AB55AAD56CB6;
defparam spx9_inst_3.INIT_RAM_34 = 288'hFC6D6608C1512D5D11A964F69B5EAEDB2B3407E9984A241288C2C35128D44A271C0E06C2;
defparam spx9_inst_3.INIT_RAM_35 = 288'hAEDF73D7EAED76BB7DDF5F277BCAD9C7536831A0409E844A2495EA34A2DDD51DA7D42C36;
defparam spx9_inst_3.INIT_RAM_36 = 288'hD389E906A85CB65F51C9646E391C8DC25ECD360AC140A050AC988D571B531DE5D3D1273D;
defparam spx9_inst_3.INIT_RAM_37 = 288'hE4122138AE56A71167945229369C56AF97CBF5FAC160BF5FAC160BE66A6CD67E57B6D6A8;
defparam spx9_inst_3.INIT_RAM_38 = 288'hD763ADD8EB75365B4DB7DBE9F4FA7E4361D0C794FA36FE8DC29E54060155325B30C69A69;
defparam spx9_inst_3.INIT_RAM_39 = 288'hD9050EC983B958AA54E9747A1F0292D5F0F97CBE16EB64AA54EA562A954AA5419FCADF2E;
defparam spx9_inst_3.INIT_RAM_3A = 288'h98D4B2773C9ED329533711982C361A8944A16130984C26130984C271B0984C2409008081;
defparam spx9_inst_3.INIT_RAM_3B = 288'hBF5F9FBB9E90AE4CA420A83864B872B1D8AB452AD990EB7EC7E433E8D3D582AF51315D0F;
defparam spx9_inst_3.INIT_RAM_3C = 288'h87D3F21B1C8DC21CCE66A30962A1512CD68C572BE65757A149A8199E5737DBEAE677BD7D;
defparam spx9_inst_3.INIT_RAM_3D = 288'h93DA755CBE5EAB97EBC65AED5CB16130560B058AF9346B3F2BD78B549A5134B36CBA9D0C;
defparam spx9_inst_3.INIT_RAM_3E = 288'hC6532994CC6EBB1B6DC7E3F2191D8ECBA5D2F972E1206517A021AE040A0D109D502B9186;
defparam spx9_inst_3.INIT_RAM_3F = 288'hD7DBB1C114A359B0F89C461F0D86BA58AA341A0D027F2E8EBEDD6EA753E9D4EA6DB71BAD;

SPX9 spx9_inst_4 (
    .DO({spx9_inst_4_dout_w[26:0],spx9_inst_4_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_4.READ_MODE = 1'b0;
defparam spx9_inst_4.WRITE_MODE = 2'b00;
defparam spx9_inst_4.BIT_WIDTH = 9;
defparam spx9_inst_4.BLK_SEL = 3'b001;
defparam spx9_inst_4.RESET_MODE = "SYNC";
defparam spx9_inst_4.INIT_RAM_00 = 288'h2709982C261A8944A16130984C26130984C271B0986C3411008081E88CD2C974B1D467D1;
defparam spx9_inst_4.INIT_RAM_01 = 288'h31304086CB7C3A5CEC349A916AC66C3A5D4F76AB055E9E4828988D67CC2A372C964F2752;
defparam spx9_inst_4.INIT_RAM_02 = 288'h66A30962B259AD188C568B3174C86C3BA2D50C165F91C7E4727ABB5DF61292EF54190662;
defparam spx9_inst_4.INIT_RAM_03 = 288'h892C05C0C16130D86C360AC13C8D46A755ECA622490EA16B35D8CC66BBA5D4FA7C399AAD;
defparam spx9_inst_4.INIT_RAM_04 = 288'hD86C3A3F209850683419ECB99E5B2618D431350A04E8894E2791E8C4FACDACF78CCAA573;
defparam spx9_inst_4.INIT_RAM_05 = 288'h8C3E1F0F86BAD8A83309FCBA3B0C7E3ADD6EB75BA9D4EA6D36DB6C95D2ED96CA65329B4D;
defparam spx9_inst_4.INIT_RAM_06 = 288'h5128944A25128944A261309C6E3511848281E88D12CB75BA58A9F2C7D3ADDF039AD9AEF8;
defparam spx9_inst_4.INIT_RAM_07 = 288'h451A8D44A251A9168B250A813E9F4828542B363361D30A8E4B255227099C4C25128944A1;
defparam spx9_inst_4.INIT_RAM_08 = 288'h7692F14EA65BB61D0ED87C566F56A3516832F8C3792E65220CC4614138C0A8DE95429EED;
defparam spx9_inst_4.INIT_RAM_09 = 288'h460A8544AF4E23522CF73AC9089D5A35DACC874BE9F70B853E5F0E66AB5186C361B1188C;
defparam spx9_inst_4.INIT_RAM_0A = 288'h4AB5A210A13C128B6EA6A2B8FE7444A311A7D50B5A173FB0DC70581BED6248F372351A8D;
defparam spx9_inst_4.INIT_RAM_0B = 288'hE8EC31F6EA6D36DB8DB75BA9B4DA6D36994CA5D32D94C864329B8ED8F4426543AA592E97;
defparam spx9_inst_4.INIT_RAM_0C = 288'h61309C70361184C281E90D16ED86C2DD2C54D85BEDFF139AD9EF197C3E231187BAD8A812;
defparam spx9_inst_4.INIT_RAM_0D = 288'h150A4522904824522A149A918CD87D42E35117119C4C25128984A15128944A25128944A2;
defparam spx9_inst_4.INIT_RAM_0E = 288'h56231DD2E56A30D9EAB3D1A4D0682B1102404148C0A6EF9E46A0EE55A2CD44A25128D46A;
defparam spx9_inst_4.INIT_RAM_0F = 288'h0763594488523AA150D96CB65D2E974BA5B2A843DDCAE56A351A6D1512F9709453315A6C;
defparam spx9_inst_4.INIT_RAM_10 = 288'hE74B05386F3C26D326C5031A1941B964B2390C7DEE9127833D5C6D260AC542A04F27920B;
defparam spx9_inst_4.INIT_RAM_11 = 288'hB6D36994DA6D36992CC6DB2992C86D3BA032E904C68765BB61B0D87B1D46931855124BA7;
defparam spx9_inst_4.INIT_RAM_12 = 288'hE9151AEF97CBE5B0B62984BE2335A359F1398C461F0F76B1D025D0B75BA9B4DA6DB71B8D;
defparam spx9_inst_4.INIT_RAM_13 = 288'h249A8D66B56BBA1F101719E04C25128984A15128944A25128944A251309C6E361184C2A2;
defparam spx9_inst_4.INIT_RAM_14 = 288'h5251B93C9B330C802041D17CC2EFA6CE60EE55AAD146A351A9148A150A85209048241209;
defparam spx9_inst_4.INIT_RAM_15 = 288'hEA753A9F4FA7D7EBF5E9ECEE5318833D5C8E252B058A7F31AA5D9025FA793A993399CCA4;
defparam spx9_inst_4.INIT_RAM_16 = 288'hD5835A1952C268F439FC7DF6B5388C41DEAE261B0960A151B0980BD603AD8484413B67F4;
defparam spx9_inst_4.INIT_RAM_17 = 288'hB6D329B4ED87C86654098D0ECB76C3E5F2F96C1D8EA34472A30B045553619E8D3222D5A9;
defparam spx9_inst_4.INIT_RAM_18 = 288'h7BA54E8945AB59EF187C35D6C74197C2DD2D96536DB8ED76BB5B8DB6D32994CA65B6994C;
defparam spx9_inst_4.INIT_RAM_19 = 288'h2721E86C35128984A15128944A25128944A25128984E351184C2A2E91D5F1198D46A32F8;
defparam spx9_inst_4.INIT_RAM_1A = 288'h51D9B4BCDFAF52A10F45A2D168A351A9148A359AC944A2492492493522D166B362B59CCE;
defparam spx9_inst_4.INIT_RAM_1B = 288'h2B0DBEBB4C9D4A22D0675C19F09D2699150DD3C15488300804440141392CD46520844040;
defparam spx9_inst_4.INIT_RAM_1C = 288'h1C8E3AD32784C2A10F573395A4B363B99C4CD5037184813E32E6570B0582C160B0582C36;
defparam spx9_inst_4.INIT_RAM_1D = 288'h2A1D52CD87CC66351A6CCE8ABF2098B00A069222B1CCCD3F9A946E17139A3740BA65347A;
defparam spx9_inst_4.INIT_RAM_1E = 288'h3B153E5D0C753616CA95DB75DF018043DFCEC6DB2994CA65B6DB4C864B6DDD1299D06813;
defparam spx9_inst_4.INIT_RAM_1F = 288'h5128944A25128944A25128944C251184C2A2F9256313A9D4EAB53A9CB5D6CB55AA552AB6;
defparam spx9_inst_4.INIT_RAM_20 = 288'h562B198AB55A2CD66B361ACD66B351A8D46A3522D588C56B39DECF37322C8E3512898481;
defparam spx9_inst_4.INIT_RAM_21 = 288'h7864A236AD238984E3B2A8D048220904C4611018504A341989048231D16894BEAFD2E34F;
defparam spx9_inst_4.INIT_RAM_22 = 288'h984C21EEE673BDDECF15F2E96CA14224A0572B960B0783C1E0F0783C15C6E16FB7576993;
defparam spx9_inst_4.INIT_RAM_23 = 288'h6D4692C12093BA92E89269D974D44E94D02ECAD522754DB0E0F2792C963ED32785472371;
defparam spx9_inst_4.INIT_RAM_24 = 288'hB6EB82052491C8E230E7E36992BA65B2992C975BFA2332A15468141A150EC976C3E6353A;
defparam spx9_inst_4.INIT_RAM_25 = 288'h5128944A24098502C209256313A9D56EF75AAD3E5AEB64A950683409F4B1F2D8642E170A;
defparam spx9_inst_4.INIT_RAM_26 = 288'h0582C564A2512492290512D18CE77CC2631037B2708E35128984815128944A25128944A2;
defparam spx9_inst_4.INIT_RAM_27 = 288'h71100806120080C040301814504A3519C88211411C6CACA752A14F8743A1B0D76331166B;
defparam spx9_inst_4.INIT_RAM_28 = 288'h76EAA552C44F9F1A384C26130984C26130982C160B0582C15C6C16DA7D6A5CC1350DC4C1;
defparam spx9_inst_4.INIT_RAM_29 = 288'h14C974F6DA669B4B0B8E1E72D55BAF5C2E380B963ED5298E4B6571C94C2615087AB99F52;
defparam spx9_inst_4.INIT_RAM_2A = 288'h0873AD92CA6532992CD87C42633098506A55098CC68764BB61F31A7E05DAEF5A73B59AC6;
defparam spx9_inst_4.INIT_RAM_2B = 288'h092D6715A9D56EF77B9DBE5AED64A8D02613F96C29D0C85CAE976BD77BC629359ACD2492;
defparam spx9_inst_4.INIT_RAM_2C = 288'h36A355CEF884C2A35158426C6E27128542E35128944A25128944A250A8582A140A050282;
defparam spx9_inst_4.INIT_RAM_2D = 288'h309850505C3E9E8AC33010144A99804B210F773B9DCEE66AB5188C048A8D46B35128540A;
defparam spx9_inst_4.INIT_RAM_2E = 288'h2C1E4F2581C0E0B0794C1E0F0782C964B0580BED82EF203B8A46C261204806030180C060;
defparam spx9_inst_4.INIT_RAM_2F = 288'h07BE9337579BCBAB93DA64EE772C9ECF2572C95CA62EF673BA5F4FA91BBD78B751A698D2;
defparam spx9_inst_4.INIT_RAM_30 = 288'hE98D0AA553B2592C5408EC29F911AB61B0B85C1D827D1B7CBA1D0EC57964849973339146;
defparam spx9_inst_4.INIT_RAM_31 = 288'h8D3E5B0B74A9D025B0A64B216EB75C2E594CE6FB8A2935AB5568B41873ADB6DA6D371FF1;
defparam spx9_inst_4.INIT_RAM_32 = 288'h6862C4D648128542C241209048241209048250A8582A140A050282F89CDEF59BDD6EB75B;
defparam spx9_inst_4.INIT_RAM_33 = 288'h30209C88867742DEEE974BA5D0E76B3558AC66331566A250A8966B46AB9DF30A8D46A331;
defparam spx9_inst_4.INIT_RAM_34 = 288'h3B9DCF0783C1E0F0783C85CB17465616C8E261204C0603010080803018504E4A359A08A2;
defparam spx9_inst_4.INIT_RAM_35 = 288'hC9E4F27B3C9E4F67B3E9ECEE530773359ACDA8B3CD9EC951A195ADEB160B0171C0E02E37;
defparam spx9_inst_4.INIT_RAM_36 = 288'hE85BDDAEEC8850AA550A05025F1D853A1CEE063230BA655D3999E8555D533B6592C6E772;
defparam spx9_inst_4.INIT_RAM_37 = 288'hA64B2170B85C2E594CC673820734A251267348F3E992CB763FE2530A1552C975BB5D6C75;
defparam spx9_inst_4.INIT_RAM_38 = 288'h41209048241209048250A8542A1409850282C80492AF88CCEA33396C3E1F0D63A7C6DF2E;
defparam spx9_inst_4.INIT_RAM_39 = 288'hB7D3A9D2E86BB598AC56231164B251AD5AEE573BE6171C95CAA331881BAD647A1B0944A2;
defparam spx9_inst_4.INIT_RAM_3A = 288'h5D16133F7D689F4B0371B0902813090080813018102C3824118481303928A4725E3ADB0D;
defparam spx9_inst_4.INIT_RAM_3B = 288'hD964AE30F569B0D64A369B099EBA52A512CA68858AFF63C2606C572B95CAE572B9E0F078;
defparam spx9_inst_4.INIT_RAM_3C = 288'hA8D46A10E76BBA5F50780B91124C33B21A29D36B87017893C663B2A9E4FA9D4D9E4B65D3;
defparam spx9_inst_4.INIT_RAM_3D = 288'h9663BE05249A4D24712873A9B6EE804866541AA596ED87C3E1AE9609641DACD76D3F21B1;
defparam spx9_inst_4.INIT_RAM_3E = 288'h50A8542A140984C281E8848EAD77C3E5F0F85BB596C53E853618EB95CAE570B85CAE572B;
defparam spx9_inst_4.INIT_RAM_3F = 288'h362359ACD773BA1F0F884C2A392C964AE552A8D451F2AE2C0D44A240A05028140A050281;

SPX9 spx9_inst_5 (
    .DO({spx9_inst_5_dout_w[26:0],spx9_inst_5_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_5.READ_MODE = 1'b0;
defparam spx9_inst_5.WRITE_MODE = 2'b00;
defparam spx9_inst_5.BIT_WIDTH = 9;
defparam spx9_inst_5.BLK_SEL = 3'b001;
defparam spx9_inst_5.RESET_MODE = "SYNC";
defparam spx9_inst_5.INIT_RAM_00 = 288'hC3491C6E36118480613018102A261A89026030C970E26F55B71B2DA753A9D2D86BB5D8CC;
defparam spx9_inst_5.INIT_RAM_01 = 288'hF50A897EAB4C259289C6650F0777CBE570F93C1DCAC150A8D8AE794C9617438179234B64;
defparam spx9_inst_5.INIT_RAM_02 = 288'hC9DCFDDC681FA196CBE3FA1A7F7B9DCA61F3C9ED3A9D4D9E4B259177BBD9C8C258A81229;
defparam spx9_inst_5.INIT_RAM_03 = 288'hD6E371FD11995068143AA59AED87CBE5F2D86B153A36F86B3198ED6743EA13098546E392;
defparam spx9_inst_5.INIT_RAM_04 = 288'h3A1D12A965BADD6CB64A94FE36F863AE170B85CAE572B95CAE572B965B79E30389C4A02F;
defparam spx9_inst_5.INIT_RAM_05 = 288'hB8DC6E572C9E4F69B4C9F52E62E3451184C240A05028140A05028140285428130984C261;
defparam spx9_inst_5.INIT_RAM_06 = 288'h301810282512890260204970C06E4DBB9F8FA7D3E9D2E974BA1D0E985432391B8D426110;
defparam spx9_inst_5.INIT_RAM_07 = 288'h64C49713ABDD6E755B5CA606BD3D9F506C782C9617458381234BE61469A8945A22888040;
defparam spx9_inst_5.INIT_RAM_08 = 288'h55C95D8F2C96C65FD2EA75369D3D9E4A610E46A30D62A048249269462B1582AE4E261288;
defparam spx9_inst_5.INIT_RAM_09 = 288'h4AA596ED87CC66753AACC5DAA52B72AD14AB77F4D6F398CADC2B72B96D2656BD2D10D38E;
defparam spx9_inst_5.INIT_RAM_0A = 288'hF8E3E5AEB75C2E554B8542E572B95CAE572B95D331BCEE77375B8C9663BE2131A0D46814;
defparam spx9_inst_5.INIT_RAM_0B = 288'hFA8DBECD185E1584C240A05028140A05028140205428130984C2616AA54A8341A150A653;
defparam spx9_inst_5.INIT_RAM_0C = 288'h304128BE5F56BFE3D2C8DC2E170B85C2E170C964B2592B8DCAE593D964AE572C9ED3EA16;
defparam spx9_inst_5.INIT_RAM_0D = 288'h7D2E06BD2C8E482A582C9E57479591A30A274579F4DC7C3308804030180C28261B8D4481;
defparam spx9_inst_5.INIT_RAM_0E = 288'hFA74F6792C9541DC8C56230D64A148A4D48A562B0D64914F2290E8549C1319CCE5EEF77B;
defparam spx9_inst_5.INIT_RAM_0F = 288'h9DCE66ED4E7B2D570D3AC67B9FEEF67171F4A964F66F074C8F0CCBB769F8FAD986C6E1B2;
defparam spx9_inst_5.INIT_RAM_10 = 288'h8542E572B95CAE572B95CAE572B95CAE170BC7FC466140A0546A55399D12AF78CCEAB79C;
defparam spx9_inst_5.INIT_RAM_11 = 288'h40A05028140A05028140205028130904C2617B2546814098CC241196C3196EB95CAE550A;
defparam spx9_inst_5.INIT_RAM_12 = 288'hE9F4F65B2C96CB65B2C9E4F2572A95CB27B4D964AE572C9F542C573C9606F54C6E9944A2;
defparam spx9_inst_5.INIT_RAM_13 = 288'h3C9E5349989A26C9E714F9FCE08C3208406130104C2A382C9608A23030987C505EC7E7D4;
defparam spx9_inst_5.INIT_RAM_14 = 288'h359ACD66A25124946A158281249448A3514854D336B5CADD6F7B3B7D2E0EBF2C8ECBEA58;
defparam spx9_inst_5.INIT_RAM_15 = 288'hBD6733B5DBEE767497C9D4B27D33789E4986B6BB3D0A8265BFA351E9ECF2571983B9586B;
defparam spx9_inst_5.INIT_RAM_16 = 288'h95C2E16EB85CB2DB8EF914CEA562B158AA14E87C466D68CCEA777C9DCEA70B4D7B321DD2;
defparam spx9_inst_5.INIT_RAM_17 = 288'h4020502813010482617BA58681309FCB5F6E75BADD70B85C2A150A85C2E172B95CAE974B;
defparam spx9_inst_5.INIT_RAM_18 = 288'hFAFD7E9D4C9DCEA753C964AE573DA7D46C576D9E87195E76994281402010080402010080;
defparam spx9_inst_5.INIT_RAM_19 = 288'hE3F1C1029B290440823090484C4A359A4AC34020503A5066CBE9D5FA7D3A9B3D9ECF67B3;
defparam spx9_inst_5.INIT_RAM_1A = 288'h2582854AA751A34F48551A564FB7D4F3BD1B6D2E12A32E8F482A584D1E4F279AA2AA49A5;
defparam spx9_inst_5.INIT_RAM_1B = 288'hEA446A4750AFB7CF455573C53C5B433362CFC96CB657177AB4D68B048A8944A148A45229;
defparam spx9_inst_5.INIT_RAM_1C = 288'h199D56EB86C2DCABB2A6DBBE2B58C3E5F53B9E4EE3094C7B36E0759D5F2BB3EBF6FAB697;
defparam spx9_inst_5.INIT_RAM_1D = 288'h6B1D429F3E963DD88A85CAE16EA54B26152B85C2E170B85CAE594C85C2DD70BA6EC06473;
defparam spx9_inst_5.INIT_RAM_1E = 288'hC9E4EE572B9ED02C572C15CAF94D6611028260A85028040205028130184C060309848261;
defparam spx9_inst_5.INIT_RAM_1F = 288'h3090080A292512068150984C584D56C4E815FA7D3E9F4FA7D3E9F4EB7D7EBB4B95CB25D3;
defparam spx9_inst_5.INIT_RAM_20 = 288'hC519DD5F8AEA6974DA6D2E4EE14E9F4FE8363C261B119FACAE8924C359B4FE7B32084041;
defparam spx9_inst_5.INIT_RAM_21 = 288'h81B2E9C09F3F36632F98C45E0CE461A914AB15128944A25124D26A159AD58CB448205069;
defparam spx9_inst_5.INIT_RAM_22 = 288'hA6C321BD05A45E6F17DCBD8EAF8ADD6DF6DACE572B95CCE776B7F6CA0D9B2DA5C8DC1F43;
defparam spx9_inst_5.INIT_RAM_23 = 288'h95C2E172B95D325B2D653AE572B85C2A554B85CB29BAFE8FC868754BBE6753A8D3E0EBF3;
defparam spx9_inst_5.INIT_RAM_24 = 288'h3C15FEB31B5E9184E240201008140A05026140984C2613098482413A04B618EA642DD50A;
defparam spx9_inst_5.INIT_RAM_25 = 288'h60984C564C564069F4FA7D3E9F4FA7D3E9F4EAF576993A9546A351C964B2592C9E4FA815;
defparam spx9_inst_5.INIT_RAM_26 = 288'h2B0D7E9D2D974C6A773B9DD2ED80AE32CB0492C1249458218442613090080A281C0D8461;
defparam spx9_inst_5.INIT_RAM_27 = 288'hA94C5E0CE46229148A15128D68B351245229048245249349A453E8943A1D22FAA0DA3054;
defparam spx9_inst_5.INIT_RAM_28 = 288'h3A255F19BEF6FB3B9D5D4EFFDFFBE3E8AF744C3EAB73B7DBEB2B8CD2C91D98EF4221A171;
defparam spx9_inst_5.INIT_RAM_29 = 288'h6542E572B85C2A152B96DBBA2533A154ECB78CCEAF95CADCE9F096D7CB5D94D089CD68D5;
defparam spx9_inst_5.INIT_RAM_2A = 288'h20180C08140A05026140A050281309848241F8E3E9B2C85BA9D52B75BADD4EA753A9D70C;
defparam spx9_inst_5.INIT_RAM_2B = 288'hE9F4FE8140A0542A15FAFD769B4C9E4AA350A8DC6E572B95CB25B3FAED2A4AFA5711C2C2;
defparam spx9_inst_5.INIT_RAM_2C = 288'h2B154AAB72B03BCD248230D86C351084406120900C28161309024060A04C544A4CBFE7B3;
defparam spx9_inst_5.INIT_RAM_2D = 288'h251A9168B3512892493522D162A253B6A170B4CA4CEC9D5CBD25EEC8DC29F2EA7E47E635;
defparam spx9_inst_5.INIT_RAM_2E = 288'hCEC6DF6BAEB5D2A9334CB6A793C8DCECF0F25430B8FAF65F9AD751C94C5DEAD4622D1469;
defparam spx9_inst_5.INIT_RAM_2F = 288'hB86C468963B158EED89D5F2F97CBE5F2B51919539548975D375DD0A7952B7DEEFF7FBFFF;
defparam spx9_inst_5.INIT_RAM_30 = 288'h40A050281409848040A6CB216EA653AA598DC763B1B4C853A9D70B854AE572B85C2E596C;
defparam spx9_inst_5.INIT_RAM_31 = 288'hFAF5369B4EA74F255187C42613098542E391A9546A2EFF599A448020100C08140A050281;
defparam spx9_inst_5.INIT_RAM_32 = 288'hA2C1186C35110440212010502A251285026150A0505449443BA5B3E9FCC28151A8D42A15;
defparam spx9_inst_5.INIT_RAM_33 = 288'h8753E9F2FD8A596E5606B270A4884F26596A76BB1D8EC86CBAE392FA05068962A9B88F84;
defparam spx9_inst_5.INIT_RAM_34 = 288'h0B962375C8DBE8AF33F619DC5E7C7227CC0EB94C19C8C35A2D1669459ACD46A3522D990D;
defparam spx9_inst_5.INIT_RAM_35 = 288'h8CD6EF95DAE572B7194AEC15648342A9D92D979DB39BEBFE7FBFDECF658623038B4A6733;
defparam spx9_inst_5.INIT_RAM_36 = 288'h85BAE14EA754B39E5139A4CE40FC6CAE150A95CAE570B85CB31DCFF98D0EA761A854EEF9;
defparam spx9_inst_5.INIT_RAM_37 = 288'h8843DDEEF773BE5F50A8D46E35057527CB0230180C06020180C28140A050281409848020;
defparam spx9_inst_5.INIT_RAM_38 = 288'h1010102A25128942A14020505649443BA5D3F98506A551B0D42A14C95CAE592E9F4F2551;
defparam spx9_inst_5.INIT_RAM_39 = 288'h79BB24DC934BA094CA66331D90C96D3A9F50C8F482454099B90FA4C35164B258230CC221;
defparam spx9_inst_5.INIT_RAM_3A = 288'h6703348E2554305089683BD5A6B25A2D568A4522D16AC66BBA9F70A8ECBE877AD670F0F2;
defparam spx9_inst_5.INIT_RAM_3B = 288'h5B74A1ACB65C329D6FC8A5AF99ECFEFFBFBD6DBCC61342CBEDF4782C161F77C8DAE46D52;
defparam spx9_inst_5.INIT_RAM_3C = 288'h5ABD5EA92F7DB214E98542E16EB7653BA0323B259AEB72B0506AB77C4EB399DBEDF2B719;
defparam spx9_inst_5.INIT_RAM_3D = 288'hA85C2A12F46E28CFA460A850060201008040301850281409844020653A9D4CA85E3864D4;
defparam spx9_inst_5.INIT_RAM_3E = 288'h402058785A4CBBE5F40A0D46A561B057A7D3A8542A372E9F536792B8D4660EF67339DD0E;
defparam spx9_inst_5.INIT_RAM_3F = 288'h56B35990CA6DBADF4F97E4363F1E91B50FA4C3596CB86C3515866110100C2A25130984C2;

SPX9 spx9_inst_6 (
    .DO({spx9_inst_6_dout_w[26:0],spx9_inst_6_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_6.READ_MODE = 1'b0;
defparam spx9_inst_6.WRITE_MODE = 2'b00;
defparam spx9_inst_6.BIT_WIDTH = 9;
defparam spx9_inst_6.BLK_SEL = 3'b001;
defparam spx9_inst_6.RESET_MODE = "SYNC";
defparam spx9_inst_6.INIT_RAM_00 = 288'hD69B99A8C259AD56AA34A29990E97D4725B3EAA62351B5C9636CF3EB94857A904CB19EAE;
defparam spx9_inst_6.INIT_RAM_01 = 288'hD915A359DEF7FF7B7C3CF58B19DFFFFFFFDE6D863EE370B75327109712ED3E581AAADA07;
defparam spx9_inst_6.INIT_RAM_02 = 288'h653AA170C97643E6753B25DF0F83AF4AE3914B462F79CCE5EEB5192A6CA5D0EA7643A213;
defparam spx9_inst_6.INIT_RAM_03 = 288'h91C8E04C150A00C06020100C261309044020653A9D4CA85EBCE6D56B3DA2CD428EB656E9;
defparam spx9_inst_6.INIT_RAM_04 = 288'h0A0D46C360AF532571974BA5F71D9F53A9B3D9E4F255197BBA1D0E87CBE5EEE366290FE5;
defparam spx9_inst_6.INIT_RAM_05 = 288'hB7EC31FB0E8B39CFA3A2D168B86D3599C64120100C2815130984A24028A09E6B4CBC27F4;
defparam spx9_inst_6.INIT_RAM_06 = 288'h34A2956ED9864FEA576DCF23879DAD53AC581C5DADE2B0563AA9327833D9CED96DBADF8F;
defparam spx9_inst_6.INIT_RAM_07 = 288'hFB05DF5DEDEDF77B9D8E65922B157ABDDECEA61A91B2981F1EDAAB34F31DCED461AD16AA;
defparam spx9_inst_6.INIT_RAM_08 = 288'h4BADDB0D71A5C19C8DD88D16ED86C3E1B0B709E469F4FC8F482855E9F4C2A987CBE5B0B8;
defparam spx9_inst_6.INIT_RAM_09 = 288'h10100C061309044020653A992C985FBD24D46BBDDECB428F3A97096542E9B8FD8FCCAA97;
defparam spx9_inst_6.INIT_RAM_0A = 288'h663B5DD10A8DCB2793D9ECF67B2B8D429F2F7743A5F0E46EAD51E5D26130943813894260;
defparam spx9_inst_6.INIT_RAM_0B = 288'hA2D168B45C351586203090080615130944815038A4806C553C27F40A8D46C36FAECEA30F;
defparam spx9_inst_6.INIT_RAM_0C = 288'hEFAEF6D960B960AE360B5539ECC355362954BA54A612EA763F5FAFE87471FB0094C251C4;
defparam spx9_inst_6.INIT_RAM_0D = 288'hAED541FEE069355ACD95BB159AB23E14938EC3529DD2E569B116A955228D46C67E4D311B;
defparam spx9_inst_6.INIT_RAM_0E = 288'h564BF65F4FA054683429FC721B1E9050AA76FA5462152C9DCF27B4DA0DAB7FEEEEF7BDBD;
defparam spx9_inst_6.INIT_RAM_0F = 288'h75429D2C9A583D24B37C35D6A7308E3A14A875D37A0322A1D92EB88CBE5B0B609CC15A8C;
defparam spx9_inst_6.INIT_RAM_10 = 288'hD9ECF2571A8CC6211098C45A0AF276AE108601F8F87A3B1C8E0703612048040201808021;
defparam spx9_inst_6.INIT_RAM_11 = 288'h20100806060C09C48030A870886D54BC25B0F98506814F9ECAE330974BA5F2FA85C767D3;
defparam spx9_inst_6.INIT_RAM_12 = 288'h0CDD820EB4532861D6CBEDF2C50A57C99810C7E3FA3D2FA7D09DE5A1C8E4744A24918682;
defparam spx9_inst_6.INIT_RAM_13 = 288'h36331D8CBF4F930B2ED87A3DA4C562AD970C642A451CA679E2B93C3C8E3EFF7EBEDB6DF7;
defparam spx9_inst_6.INIT_RAM_14 = 288'hB7E43A4355BB5D2C34095BE1D4FE8F4B6592EA159F39CFF77B3B3C2C6D5E06D35AA954AA;
defparam spx9_inst_6.INIT_RAM_15 = 288'h499C92270F6CA9D4EBE904C29F40A2DA71786CC6A36B94C15AE28D252AE5B4E86B321B8F;
defparam spx9_inst_6.INIT_RAM_16 = 288'hB95CAA4F1376ADD06512013C9A4D261309A59240D82A150A0440006532994C9655301E91;
defparam spx9_inst_6.INIT_RAM_17 = 288'h4130B0846A4BBBA3D1E9FCFE7F3E9E4AE351A7D3E5F2F985472593C95CAE571A8D46A351;
defparam spx9_inst_6.INIT_RAM_18 = 288'hBBFE4A207400B3E30DE8F4866342B25EA54AC250E06E261B0D04612010080606140DC481;
defparam spx9_inst_6.INIT_RAM_19 = 288'hB7BB38AAF35BB258CB958A392EF4BCEDB4592C863EFF7EBEDBADF70C5D4A36D964B39EB2;
defparam spx9_inst_6.INIT_RAM_1A = 288'hC84395B0FD8FCC28340A159B15BCE5F234B9FADCD9E6C35AAD548A562B156CB45DA44DA6;
defparam spx9_inst_6.INIT_RAM_1B = 288'hF99552C762AA59F1189D5F2F95C9DBE3E6EE24924D269251ADDD90F97CC28977CBE12C34;
defparam spx9_inst_6.INIT_RAM_1C = 288'h1201387A3C26938BE5E2E930963A1B89022055329D4EA753AA574CB6DB6D92B54A2659F0;
defparam spx9_inst_6.INIT_RAM_1D = 288'hD9ECFA7D3D9E4AE572C8DC2A130984C2A351A8D466351A8DC6E592DA753695247EAD8E45;
defparam spx9_inst_6.INIT_RAM_1E = 288'hE9FD0AC562B2DFE84EF3612048130984C24120904826161D1289036140F08055393763F2;
defparam spx9_inst_6.INIT_RAM_1F = 288'h463BBE719BE3E86FD62C863EE17FBF5FEE18FBF59E7CFA6C37A0F449BB4C6C340BA0690E;
defparam spx9_inst_6.INIT_RAM_20 = 288'hC8DC6E3B2E9F4F2752C8C3D5A6B45AAD168B56AAD56CB6623213221553850C867A2D96A9;
defparam spx9_inst_6.INIT_RAM_21 = 288'hADDF2FB7CCE5E92DB1A6BAD94CA764BF64352A8D46C987CB60ADD3C8D425F70D97CC2835;
defparam spx9_inst_6.INIT_RAM_22 = 288'hE2F138BE5F369689035532994CA64AA51088652A51269453B7E4D60AA5DAE750A050ECD8;
defparam spx9_inst_6.INIT_RAM_23 = 288'hE96CAE33088442213088442211098546E372D9F53A97347E2D8E4512013C9A3C1E0F0783;
defparam spx9_inst_6.INIT_RAM_24 = 288'h3479A46A130984C24120904826271D970D6571C0ECBA5036AEE3F2E9F4FA7D3E9F4F67B3;
defparam spx9_inst_6.INIT_RAM_25 = 288'h3C8E030380C7DC3038EB75A2630D7D3ADFF1D429002C32098059F2EA854EE571B1DFA88F;
defparam spx9_inst_6.INIT_RAM_26 = 288'h97BB5588C563355A8D66AB21AEC352305886723B39F6416AB4112C88AE3BB5C4C9606E16;
defparam spx9_inst_6.INIT_RAM_27 = 288'hA6BADD52CB7ECBAA164B9DCAE785C25C2B92E974FE6141A053E9F4D8D3D9CAD674BE6130;
defparam spx9_inst_6.INIT_RAM_28 = 288'h4522512A964B2592A964A2112ECB784CAA972BA5D2BF2A7D402AD8ADD72B93BAE5EDEE34;
defparam spx9_inst_6.INIT_RAM_29 = 288'h87BBDDEEF884426130A8DCB2531376298E65128944A2502F9389A3C1E0F49E51309C0DE6;
defparam spx9_inst_6.INIT_RAM_2A = 288'h20904826151C92CB457140E8944D2DAE63F3FA7D3E9F4FA7D3E815FA74F2551984421F0F;
defparam spx9_inst_6.INIT_RAM_2B = 288'hDB6DA269228CBB910610A910600C36B622970B0D92E972B15B666E4409B0903612890261;
defparam spx9_inst_6.INIT_RAM_2C = 288'hA843EE16F56AB59C2DB279D54EB23BC25E938DD71F617FBA6572582C8E030381C05C3038;
defparam spx9_inst_6.INIT_RAM_2D = 288'h5BA5CAE573B95829B2D90512CB74B0D7E9B3D8DBDDAED8753EE171A7CBE1D0F97CC26110;
defparam spx9_inst_6.INIT_RAM_2E = 288'h4432A5B90F98D4AC364B9D7E50D352B3A4D78D572B93CADD69AC138632D952CC874FEC17;
defparam spx9_inst_6.INIT_RAM_2F = 288'h67BBDDECF16629CE853321990E8642A10E46D1E0EC784F28988E6744A25128954B2994C9;
defparam spx9_inst_6.INIT_RAM_30 = 288'h60B8A4925C352E65F41A8D46A351A8D46A350AFD367719843E1F0F77BBDDEEF77BBD9CEE;
defparam spx9_inst_6.INIT_RAM_31 = 288'h41208C42108777A9F41B0D4AA552A8D6E40C23797094381B89426120984824030B0986C2;
defparam spx9_inst_6.INIT_RAM_32 = 288'h06C0A89CF2463337186D0E3AC385CAE4F0781C0602E180C7DFEE180C162EC1066598C642;
defparam spx9_inst_6.INIT_RAM_33 = 288'hF99556EB73B057675297CBE9F70C86472371E9ECF67D3E9F53A9B30A6CB6614E9E4AE310;
defparam spx9_inst_6.INIT_RAM_34 = 288'h2B7CE9CAA141261BF24BC66F77AACBDC676F96C2DD72DB7EC86AB82A8D3E9D3D9F4B63B1;
defparam spx9_inst_6.INIT_RAM_35 = 288'h53B22534AB5D2A12E9330170743B1F100A4544AA594CA652A512694553BE413E9FD0ACB7;
defparam spx9_inst_6.INIT_RAM_36 = 288'h1A8D46A351A8D42A150AFD367719843E1D0E7743A1CEF773399AAD46A34DA4CF5DA5CEA5;
defparam spx9_inst_6.INIT_RAM_37 = 288'h4A84FE5F209FCE218AD258E450281309024020100804020205428150B0A0925D3DB6A615;
defparam spx9_inst_6.INIT_RAM_38 = 288'hBA6542EB96D260B0792C8E070381C05FEE181CF60A2296208442C330905C94514140CE0D;
defparam spx9_inst_6.INIT_RAM_39 = 288'hD8F4826331A0502A151B0582C161B0D82C161B0D82C364B95BA9B3FA29FCA48861A42E58;
defparam spx9_inst_6.INIT_RAM_3A = 288'hC80CD2A95298471D0B75BA994CB55B36A012D8EC6E10F7743ADFB01A9D92E761A857A792;
defparam spx9_inst_6.INIT_RAM_3B = 288'hA4A9F89439158F880454B2594CA4522956CC97F486A350A9596EF71AFCF216D85AA954CC;
defparam spx9_inst_6.INIT_RAM_3C = 288'h0AFD3275187C39DCED7743A1D0F87BB99AAC4612C57EAE55A20CA564422556BB5DAE550A;
defparam spx9_inst_6.INIT_RAM_3D = 288'h9140582C160A84C02010100C0403030582C15030A0926E463AE8151A8D4AA551A85429F4;
defparam spx9_inst_6.INIT_RAM_3E = 288'h4C964B2792C8E07038DC0470E0131390C4006110102A20071AC74A8B14FA3D1F97499F29;
defparam spx9_inst_6.INIT_RAM_3F = 288'h1C8E070381C0DC6C16DAA60B1F73C1E06C5709FCDD323354B74F56EA8DC6FB5EAAE5F499;

SPX9 spx9_inst_7 (
    .DO({spx9_inst_7_dout_w[26:0],spx9_inst_7_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_7.READ_MODE = 1'b0;
defparam spx9_inst_7.WRITE_MODE = 2'b00;
defparam spx9_inst_7.BIT_WIDTH = 9;
defparam spx9_inst_7.BLK_SEL = 3'b001;
defparam spx9_inst_7.RESET_MODE = "SYNC";
defparam spx9_inst_7.INIT_RAM_00 = 288'h95D2E970B451A9996EC863E5EED563B71DF00A0D46BF4FA9592C76F984C27F3E9F502C57;
defparam spx9_inst_7.INIT_RAM_01 = 288'h64B25526934AAE9DB0FA7D3ABF64BC61AC745BA5526B338E359469454B6DD2D7642E14E9;
defparam spx9_inst_7.INIT_RAM_02 = 288'h67339DF0F77234D86C360AF958AC552610A683C1E1108955AED76B953200B2291693C9A3;
defparam spx9_inst_7.INIT_RAM_03 = 288'h20100402020A09C92561A89C724F3FBF6DF73A9546A150A8D46A35FA6CEA31077BB9DAED;
defparam spx9_inst_7.INIT_RAM_04 = 288'h0420C84228298801AEAB0A8012242CA38A8B1AFCC2412090CA5F8991B89C4A120100C240;
defparam spx9_inst_7.INIT_RAM_05 = 288'h098D42C374CBE974590BAE5E246F2AA4D5C9E7F5F2C171BBCB28575D8E4F4BB1C8E47396;
defparam spx9_inst_7.INIT_RAM_06 = 288'hA5CAD946945C3B63F209642E1F45BBE4EDD41A150A632F974FA9F6EB16130370B0DBEB94;
defparam spx9_inst_7.INIT_RAM_07 = 288'hEA8D92C952B15DB15A5D46E74F84B1539D0945AADD50984BA594CA85BADD6EB6522914AA;
defparam spx9_inst_7.INIT_RAM_08 = 288'h358AFD58AA4C21CEC7632998F29B55AA53097411F4923A1E12C72253B2594AC77547A9F5;
defparam spx9_inst_7.INIT_RAM_09 = 288'h61A8944E3D373B2A171A053E7F40A0D46814F9ECAA31087C3A1D0D773B9DCCE56A34D84C;
defparam spx9_inst_7.INIT_RAM_0A = 288'h9A432076A4A64306070A74FE433299D3220CD2C0982C24018102403018080413128E4B66;
defparam spx9_inst_7.INIT_RAM_0B = 288'h5C8DDA2E9E29A157C8C36999630BA9602D53AADDBAE595D8E7E10410A0B0E621098585EE;
defparam spx9_inst_7.INIT_RAM_0C = 288'hB7E47A6352B1DCEC764A84ADEEC76CBF6615DA7542A162B9DD2E776BADD2E773B9DD32B9;
defparam spx9_inst_7.INIT_RAM_0D = 288'hCEEF737397C358212B3522952A874C2E9B6ED7DBA5B0C45124D2AA85C2D9469353B69F4F;
defparam spx9_inst_7.INIT_RAM_0E = 288'h8431D8F29B54214EA633712C784E2E1246C1443AE9B6FE9050AC564B95427F20A1DA337B;
defparam spx9_inst_7.INIT_RAM_0F = 288'hE9ECB65D30A053E7D2D8DC21EEF87C3A1CED66AB55A8D46A31188C2512815A9A441DCF07;
defparam spx9_inst_7.INIT_RAM_10 = 288'hEDBDC69B2D90D0293133C8942E250980C04020100804130A8E094571A090281A253267D6;
defparam spx9_inst_7.INIT_RAM_11 = 288'hE400082C3B2E3925759A860F5F8499A9040072000000020D1142E254591D2546A1489A4F;
defparam spx9_inst_7.INIT_RAM_12 = 288'hD8539D6CA75C365F30B854324155C3E6335A9CBE17077FA64FA8986CFFBEA67F2F178D2C;
defparam spx9_inst_7.INIT_RAM_13 = 288'h351A51289654B76012298CBA14E458A452AA663B1D6AA452AD58CC875C428763B9D8AA54;
defparam spx9_inst_7.INIT_RAM_14 = 288'h32F93C8664381AC923454B7A2544AAD92C551AEC69D6E092DA333ACE5EEB539ACC5C230B;
defparam spx9_inst_7.INIT_RAM_15 = 288'hC853E5F2FB853E1CCD56B355A8C46235186C150A815C9C45A29127A4BA18F08742190AC6;
defparam spx9_inst_7.INIT_RAM_16 = 288'hC5E9140E160984802010100804020A09C72461204C28181B292333D8E4723B2F9FCFA591;
defparam spx9_inst_7.INIT_RAM_17 = 288'h3975F2DAFE3904434541081154C92000414302C07161466EC3E79388442E3F30A1542B32;
defparam spx9_inst_7.INIT_RAM_18 = 288'h86BB69E348C4E6B59B9D3612E56D93BE63F5BDFFBEBE5E289FCCA93510484821098A8B0C;
defparam spx9_inst_7.INIT_RAM_19 = 288'h5B2D4E9D186928928A663B21AEC65AA914AB97EC86A975B9D7A32E65BAE174BA642D966A;
defparam spx9_inst_7.INIT_RAM_1A = 288'h675C468B66BAD86BD377AB5574D28BDA30F99D4EAB559AC3D79EAA552A996EC96E43E434;
defparam spx9_inst_7.INIT_RAM_1B = 288'h97CBE1ECE67339184B057A793E9F4F26D1277431DD108639950AE6431954D28740970984;
defparam spx9_inst_7.INIT_RAM_1C = 288'h2090482412018544E35098502C2A22A45CB0B85C321B1E8F472370C864321B1E8EC69EEE;
defparam spx9_inst_7.INIT_RAM_1D = 288'h00412EA583420150F1E611C4E4EC89D2A1B3262BB22340A053E95247A1E8523712850261;
defparam spx9_inst_7.INIT_RAM_1E = 288'hBDBE5B0D71A5C6E3F45C15DB2D1713050FE565925048292188848272022CC000028D0441;
defparam spx9_inst_7.INIT_RAM_1F = 288'h35AADD90C7632DD90CE90D0EC5509EC65AAB85CAE570A74AA5548A54AAA5A539C566F59B;
defparam spx9_inst_7.INIT_RAM_20 = 288'h6723116EBD71CDED19BDE6EF5185A8465889553B29DB0E97CC28345BADDAC74C82B114AA;
defparam spx9_inst_7.INIT_RAM_21 = 288'h167AF95EAF5726D107744A7156A84A9CCA653329A0F28638974784A8FD0ECB74B957A751;
defparam spx9_inst_7.INIT_RAM_22 = 288'h50A060564E2B27DA4E76C3A9F90C86472391C8E4763D1D8DC25EEE97D42A10F985C25ECE;
defparam spx9_inst_7.INIT_RAM_23 = 288'hA942B1BF6F9FCAA1F3298CCA613D8ECBE9D3885284BC5A240DC6A320900402010100C0A1;
defparam spx9_inst_7.INIT_RAM_24 = 288'h0B6D6F93BA5C8B89C354EBA060030B0E484261B9186A36198882A371A04D14B13EB0AC77;
defparam spx9_inst_7.INIT_RAM_25 = 288'h0AADDADF276AAD56CB85CAE972A65225148A44AAA58116ACE2B57BEEDEEB5386B1506876;
defparam spx9_inst_7.INIT_RAM_26 = 288'h4A9D469D1A6BAD54AA554B7A2543B1D8AC352B9D92C74E843556CA149A954CB663325B8F;
defparam spx9_inst_7.INIT_RAM_27 = 288'hD57AFD9ABD5EAE5286544A6D569943A10E47FA1592E973B95BEBB3D9CC0D8082443022B5;
defparam spx9_inst_7.INIT_RAM_28 = 288'h152321D4FA7DC365F3E974BE5B1B8D421F0F985426110A86CB653067A38980BE56A69127;
defparam spx9_inst_7.INIT_RAM_29 = 288'h974BB6032F8F47633077EAD9046D2D1648C32090480402018140C181B8AC9C5F299E556A;
defparam spx9_inst_7.INIT_RAM_2A = 288'hF2C2D13032020986415198906C331084C4837118205027083674971A1BF6AF96753FA1D1;
defparam spx9_inst_7.INIT_RAM_2B = 288'h34AAA174CA6431D8AC65C2E596EF8ADA355BCE5EE72D63A150EC989D2642E796D4CE5245;
defparam spx9_inst_7.INIT_RAM_2C = 288'h765BFE6975C260EC551B05429D2B7BB196EB5522554AB55AB25DB10B25D2B8F4512514AA;
defparam spx9_inst_7.INIT_RAM_2D = 288'hB67341A0C169B85DACFA1592E984C2E170775C056202AE389D976E85BB1D8AB449A514CB;
defparam spx9_inst_7.INIT_RAM_2E = 288'h2A954A9F3C8D42E391D96CAA2EF7854660CEA94C59E4CE55A69148F5833D9AB06B40DDAB;
defparam spx9_inst_7.INIT_RAM_2F = 288'h376AE5287E2D964AA36130984C260B8A4543B25134BE6E27950EA7C3829990E97DC3E655;
defparam spx9_inst_7.INIT_RAM_30 = 288'h41B910400E45D9E8E450E11D4E9E2E30EE15A7CC05DEC87659E67218E3EDD8FB7DBF212F;
defparam spx9_inst_7.INIT_RAM_31 = 288'hA763A9B0CA70D1B11B7D3E92FF3B86C42A582BA65F69A1C2E4ECEF8509A54073020502E3;
defparam spx9_inst_7.INIT_RAM_32 = 288'h1B753255076AAD970BA5C2DD6CA351ADDD91FB0DBE54E75BA952282492512EBA6E3F6190;
defparam spx9_inst_7.INIT_RAM_33 = 288'hE9854EE986CC6A773B9DAE7EB2F4511C9049542A5D50B8532956ACA76C068975CA60EC56;
defparam spx9_inst_7.INIT_RAM_34 = 288'hD9DC6E391B8C3D184B56AB61F10471345BEB1672B158AF6A4060ECD7F3D9649E744C1E88;
defparam spx9_inst_7.INIT_RAM_35 = 288'hC2D928743B26170B65A27178962B09120D47D49319A8C25232DFF2F99512A54F9F4B6592;
defparam spx9_inst_7.INIT_RAM_36 = 288'h53ECCEE7024616233056DBCE6F57A2D12895F963F1F90B85C6E2EFE5D2652A802F940DE5;
defparam spx9_inst_7.INIT_RAM_37 = 288'h287BEDD2DA7EC428551A1D8EE783C15FE951D9525110C8280143226140CC422C3EBF1BE6;
defparam spx9_inst_7.INIT_RAM_38 = 288'hB6CB65D4E95B29DD930A6CA5CCB65431D8AC64F1C557109A55AC54FA74ADF2CA5F341E10;
defparam spx9_inst_7.INIT_RAM_39 = 288'h5D2E52E13768A0D12A364BF2391A83395B2EC87C8AA763B25CEC56F953D58CB85BADD6EB;
defparam spx9_inst_7.INIT_RAM_3A = 288'h3602C182C061BE6352377B05A4EF6DB29AEC14C9608AAB689D84E2E7B36A4F9AE46A355C;
defparam spx9_inst_7.INIT_RAM_3B = 288'hA1E934962E1B9F964C469B05609E47211990B87C8E833F96CB65B2983BE1F3097CBE1C8C;
defparam spx9_inst_7.INIT_RAM_3C = 288'h97E4064935A2D128955A7C761D1F904FA50EF5C214EA753AA0CFC4037978BA4D2E170944;
defparam spx9_inst_7.INIT_RAM_3D = 288'hD874BE8363C25C29B28733951C603E1644A0815120821315978B637825A3394E6C4AF40B;
defparam spx9_inst_7.INIT_RAM_3E = 288'hD9D459A6A44BAE18EC865BD2DBBFEFF2B4976C0521C69443A616EBA653218EC86CBAA191;
defparam spx9_inst_7.INIT_RAM_3F = 288'h98647E7F3B8C3EE0121A1D4EC562B15869F3C84B9D92CA6532994C75AAD58EC9542E9DD3;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[30:0],sp_inst_8_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b00;
defparam sp_inst_8.BIT_WIDTH = 1;
defparam sp_inst_8.BLK_SEL = 3'b000;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFFFFFF211FFF3FFFCC003F7C4023FFE03FFFE07FFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_01 = 256'hFFF07FFFE0FFFFFFFFFFFFFFFFFFC4E0FF8FFFCC001FFE3023FFF03FFFE0FFFF;
defparam sp_inst_8.INIT_RAM_02 = 256'h7FC40003FFEC23FF80783CE3FFFFFFFFFFFFFFFFFF300E7FE3FFC4000FFEF823;
defparam sp_inst_8.INIT_RAM_03 = 256'hFFFFFFFDC30FFE1E640003FFF623FF000000F7FFFFFFFFFFFFFFFFFFE6301FF8;
defparam sp_inst_8.INIT_RAM_04 = 256'h7FFFFFFFFFFFFFFFFFFFFF24C3FF86040000EFD333FF0000007FFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_05 = 256'h7FE7F1FE0000007FFFFFFFFFFFFFFFFFFFFFE921FFF8060000FFCB33FE000000;
defparam sp_inst_8.INIT_RAM_06 = 256'hFF6C3FFF12000E1FF1B9FC0000003FFFFFFFFEFFFFFFFFFFFFFD01FFF8060001;
defparam sp_inst_8.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFD99FFFFF000F0FFBF9FC0001803FFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_08 = 256'h000F003FFFFFFFFFFFFFFFFF07FFFFF283D9FF000F47F9FCFC0007803FFFFFFF;
defparam sp_inst_8.INIT_RAM_09 = 256'h3F800FC3FCF8FF800F003FF380FFFFFFFFFFFF27FFFFFCE7F1FF800FC7FD78FF;
defparam sp_inst_8.INIT_RAM_0A = 256'hCFFEFFFFFFD9F00FC00FC0FE78FFC00701FFFF00FFFFFFFFFFEF0FFFFFFF27E0;
defparam sp_inst_8.INIT_RAM_0B = 256'h3F007FFFFFFFFFC7E0FFFFFFF6F807C01FC07F7C7FE00003CD7F007FFFFFFFFF;
defparam sp_inst_8.INIT_RAM_0C = 256'h16FE7FF00000003F807FFFFFF79FFBC0FFFFFFFD7827C03FC0337C7FE0000383;
defparam sp_inst_8.INIT_RAM_0D = 256'hFF0FAE06DDFFC01FFE7FF00000007F80FFFFFFFF713FE0FFFFFF8F5C016FFFC0;
defparam sp_inst_8.INIT_RAM_0E = 256'hFFB986C837FFFFF803EB0FEFFFC00FFEBFF8000000FFC1FFFFFFDC421D38FFFF;
defparam sp_inst_8.INIT_RAM_0F = 256'hF001001FFFFFC7FFFA0E1018FFFFE021F78FEFFFE007FF3FFFE00000FFE7FFFF;
defparam sp_inst_8.INIT_RAM_10 = 256'h0FFFE0023FB7FFF833800FFFFFEFFFFE19600FFFFFC0E0FBE39FFFE0067F3FFF;
defparam sp_inst_8.INIT_RAM_11 = 256'h1D7FF003FFDF7107FFF0011FC7FFFE030000FFFFFFFFFE3FC023FFF801F97CE2;
defparam sp_inst_8.INIT_RAM_12 = 256'h3E0FFFFFFF0030163C000FFFF3B83BFFF800CFC3FFFF0700007E07FFFFFFBE00;
defparam sp_inst_8.INIT_RAM_13 = 256'h63E7FFFF8000000E03FFFFFF00472DF0001FFFFF5C39FFFE00CFE7FFFF000000;
defparam sp_inst_8.INIT_RAM_14 = 256'hFFFFF728EFFE0163F7FFFFC0F000040003FFFF803CF900001FFFFF8E11EFFE01;
defparam sp_inst_8.INIT_RAM_15 = 256'h7FC01F8E00003FFFFF6B947FFE81F3F7FFFFC7F8000000000FFFC0003F00001F;
defparam sp_inst_8.INIT_RAM_16 = 256'h1E3800000000001FC0007C30013FFFFFB5CC7FFF03FFD7FEFF8F380000000000;
defparam sp_inst_8.INIT_RAM_17 = 256'h7FFFFFFFFBFFF83C380000000000078000000001FF0FFFFEC2FFFF87FFDBFE3C;
defparam sp_inst_8.INIT_RAM_18 = 256'h0000FC3FFFFEB0FFFFFFFFF5FFF9F8F80000000000030000000000FF07FF6D60;
defparam sp_inst_8.INIT_RAM_19 = 256'h00000000800000000379FFFFFFD83FFFFFFFFE1FF1F0FE7CC000000001800000;
defparam sp_inst_8.INIT_RAM_1A = 256'hFF03F9FFF7C03CC0000000800000000371FFFFFFE89FFFFFFFFF03F1E1FBF731;
defparam sp_inst_8.INIT_RAM_1B = 256'hF03FF40FFFFFFFFF03F9FFEF0FF7C0030000800000000683FFF8FFBC1FFFFFFF;
defparam sp_inst_8.INIT_RAM_1C = 256'h8000001F0007FF803F7B07FFFFFFFFC1F8FF1E3FFA610700008000000F0003FF;
defparam sp_inst_8.INIT_RAM_1D = 256'h3CFFFE200780008000003F80FFFF003FB197FFFEFFFFC070FEBEFFFC21078000;
defparam sp_inst_8.INIT_RAM_1E = 256'h7FFFCCFF60000039FFF8310300000000007F0FFFFE0000B0CB7FFE3FFFE0007C;
defparam sp_inst_8.INIT_RAM_1F = 256'h1FFFE000000071FBFFF03FF0000001FFEC000108004000007F0FFFF800004163;
defparam sp_inst_8.INIT_RAM_20 = 256'h0018004000007E0FFF8000000FA2FFC0001FF000003EFF90200018004000007E;
defparam sp_inst_8.INIT_RAM_21 = 256'h7800003FFE00200000004000007F0FFF0000003FD9CF87800EF800003FC0C020;
defparam sp_inst_8.INIT_RAM_22 = 256'h03FFF4E78F0000B80000178000000000004000007FDFFE0000017FE8E78F8006;
defparam sp_inst_8.INIT_RAM_23 = 256'h00007FFFC00C000FFFEB720FC000BDFFC0130000100000004000007FFFF80000;
defparam sp_inst_8.INIT_RAM_24 = 256'h000010000000400000FFFF803F001FFFFB3A07C0007DFFF01000001000000040;
defparam sp_inst_8.INIT_RAM_25 = 256'h6000003EFFFFA8000014000000400000FFFF003F803FFFF199C3C0007BFFFF18;
defparam sp_inst_8.INIT_RAM_26 = 256'h003F81FF07E04EA000001F7FFFE80000100000006000007FFE003F807F8FE09C;
defparam sp_inst_8.INIT_RAM_27 = 256'h00001000007FF0001F87FF8000277000001F6FFFEC0000100000003000007FF8;
defparam sp_inst_8.INIT_RAM_28 = 256'hBFE3F4800018000000080000FFC0001F0FFFC000230000009FBFFFF400001800;
defparam sp_inst_8.INIT_RAM_29 = 256'hF0FE0990000007BFE3F5800008000001480000FF0000001FFFF03E13A000000F;
defparam sp_inst_8.INIT_RAM_2A = 256'h00F80000007F3FF0FF04D0000003DFE1F4900000000003E80000FF0000003FFF;
defparam sp_inst_8.INIT_RAM_2B = 256'h000B000003E80000E0000003FE1FF1FF1CE8000003DFF3F4300000000003E800;
defparam sp_inst_8.INIT_RAM_2C = 256'h000001E7C3FC00000A000001C80000C0000003FE0FFFFE7C74000000EFF1F400;
defparam sp_inst_8.INIT_RAM_2D = 256'h3FFF807FF0FE9A000000FA01F80000081F00000800000000001FFF0FFFFEFD34;
defparam sp_inst_8.INIT_RAM_2E = 256'h0004000001F0007FFF807F80FECC0000075C007A0000083F00000C0000000000;
defparam sp_inst_8.INIT_RAM_2F = 256'h0002000008FC000006000003F001FFFF807F8FFE0F00001E4C003A0000087F00;
defparam sp_inst_8.INIT_RAM_30 = 256'h7F8013C001F1BC000200000AF8000006000003F801F8FF817FBFD82780007C2C;
defparam sp_inst_8.INIT_RAM_31 = 256'h07F81FF80787007F901B4003CFBC000A00001AF0000006000003F803F87F833F;
defparam sp_inst_8.INIT_RAM_32 = 256'h1800000007C00003F06FFC001F807F8009A017C09C090000001A700000078000;
defparam sp_inst_8.INIT_RAM_33 = 256'h1ED11E463C00001800000007C00000007FFC003F03FF0006C02FC09E103D0000;
defparam sp_inst_8.INIT_RAM_34 = 256'h01FE1C000001607FFB0F007C80000C00000007C0000001FFFE01FE03000002F0;
defparam sp_inst_8.INIT_RAM_35 = 256'h07FF070007C1FF01FE7C00000039F7FF0405FCC0000401000007F80E0007E3FF;
defparam sp_inst_8.INIT_RAM_36 = 256'hC9000005FF80000FFFC3001380FE03C07C0000901FDFF9C804FC800004FF8000;
defparam sp_inst_8.INIT_RAM_37 = 256'hFF6FAC67FF0001C1000005FE80001FFFC1003F807C0100FC3FFFFC5F3FFD900A;
defparam sp_inst_8.INIT_RAM_38 = 256'h7FFC0000008EF07CFFD699FE814DBD000004FF00003FFFE0000FF8000000E763;
defparam sp_inst_8.INIT_RAM_39 = 256'h0C00001FFF8007EFFE0000001FC13FFFD6261E01599C000005CF00003FFFC000;
defparam sp_inst_8.INIT_RAM_3A = 256'h1030B00E8000040000001FFF9C1F8FFE01C0003F001FF1D1046400BCE6800004;
defparam sp_inst_8.INIT_RAM_3B = 256'h0078001FF8E2C0401AE41C4000040000007FFFFC3E0FFC01E0003C001FF0C581;
defparam sp_inst_8.INIT_RAM_3C = 256'hFFFF7C03E01FF000E0001FFFB8C0003F60F06000060000007FFFFC3C07FC03F0;
defparam sp_inst_8.INIT_RAM_3D = 256'h70000381E0000FB1C17FC8001FE000E00007FFFB60000390107000070000000F;
defparam sp_inst_8.INIT_RAM_3E = 256'h83FC7006A83F00FA00078070000179F97FC0003F8000400007E3FEF000371780;
defparam sp_inst_8.INIT_RAM_3F = 256'h01FE0000003FC0001E28006A3F84FE80060C3000004F9C1FF0003F0000804F03;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[30:0],sp_inst_9_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b00;
defparam sp_inst_9.BIT_WIDTH = 1;
defparam sp_inst_9.BLK_SEL = 3'b000;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'h00000000000000000000FFFFF0000080001FFFFFC0001F800000000000000000;
defparam sp_inst_9.INIT_RAM_01 = 256'hFFFF80001F0000000000000000000000007FFFF0000000001FFFFFC0001F0000;
defparam sp_inst_9.INIT_RAM_02 = 256'hFFF8000000001FFFFF87C31C000000000000000000C000001FFFF8000000001F;
defparam sp_inst_9.INIT_RAM_03 = 256'h000000FE000001FFF8000000001FFFFFFFFF08000000000000000000F8000007;
defparam sp_inst_9.INIT_RAM_04 = 256'h80000000000000000000FFC000007FF8000010200FFFFFFFFF80000000000000;
defparam sp_inst_9.INIT_RAM_05 = 256'h00180FFFFFFFFF80000000000000000000FFF0000007F8000000300FFFFFFFFF;
defparam sp_inst_9.INIT_RAM_06 = 256'hFF800000EC0000000C07FFFFFFFFC0000000000000000000FFFE000007F80000;
defparam sp_inst_9.INIT_RAM_07 = 256'h000000000000FFFFE00000000000000407FFFFFFFFC0000000000000000000FF;
defparam sp_inst_9.INIT_RAM_08 = 256'hFFFFFFC00000000000000000F8FFFFFC0000000000000603FFFFFFFFC0000000;
defparam sp_inst_9.INIT_RAM_09 = 256'h000000000307FFFFFFFFC00C7F000000000000F8FFFFFF0000000000000207FF;
defparam sp_inst_9.INIT_RAM_0A = 256'h3000FFFFFFE000000000000187FFFFFFFE0000FF000000000010F0FFFFFFC000;
defparam sp_inst_9.INIT_RAM_0B = 256'hC0FF80000000003800FFFFFFF800000000000083FFFFFFFC3280FF8000000000;
defparam sp_inst_9.INIT_RAM_0C = 256'h0901FFFFFFFFFFC07F80000000000400FFFFFFFE00000000000C83FFFFFFFC7C;
defparam sp_inst_9.INIT_RAM_0D = 256'hFFFFC0000000000001FFFFFFFFFF807F000000000EC000FFFFFFFF8000000000;
defparam sp_inst_9.INIT_RAM_0E = 256'h000079F008FFFFFFFFF0000000000001FFFFFFFFFF003E000000003DE000FFFF;
defparam sp_inst_9.INIT_RAM_0F = 256'hFFFFFFE00000380001F1E007FFFFFFFFF8000000000000FFFFFFFFFF00180000;
defparam sp_inst_9.INIT_RAM_10 = 256'hF0000001C07FFFFFFFFFF00000100001E08000FFFFFFFFFC006000000180FFFF;
defparam sp_inst_9.INIT_RAM_11 = 256'h3EFFFFFFFFFF80F8000000E03FFFFFFFFFFF0000000001C0001CFFFFFFFFFF01;
defparam sp_inst_9.INIT_RAM_12 = 256'hC1F0000000000039FFFFFFFFFFC0FC000000303FFFFFFFFFFF81F80000000000;
defparam sp_inst_9.INIT_RAM_13 = 256'h1C1FFFFFFFFFFFF1FC000000003810FFFFFFFFFFE07E000000301FFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_14 = 256'hFFFFF81F1000001C0FFFFFFF0FFFFBFFFC0000001F00FFFFFFFFFFF03E100000;
defparam sp_inst_9.INIT_RAM_15 = 256'h80000070FFFFFFFFFFFC0F8000000C0FFFFFF807FFFFFFFFF000001FC0FFFFFF;
defparam sp_inst_9.INIT_RAM_16 = 256'hE007FFFFFFFFFFE0000000FFFFFFFFFFFE07800000000FFFFFF007FFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_17 = 256'h8000000007FFFFC007FFFFFFFFFFF8000000FFFFFFFFFFFF070000000007FFFF;
defparam sp_inst_9.INIT_RAM_18 = 256'hFFFFFFFFFFFFC18000000003FFFE0007FFFFFFFFFFFC000000FFFFFFFFFFFF83;
defparam sp_inst_9.INIT_RAM_19 = 256'hFFFFFFFF000000FFFFFFFFFFFFE0C000000001FFFE0001FF3FFFFFFFFE000000;
defparam sp_inst_9.INIT_RAM_1A = 256'h00FFFE000FFFC33FFFFFFF000000FFFFFFFFFFFFF06000000000FFFE0007F80E;
defparam sp_inst_9.INIT_RAM_1B = 256'hFFFFF83000000000FFFE001FFFF83FFFFFFF000000FFFFFFFFFFFFF060000000;
defparam sp_inst_9.INIT_RAM_1C = 256'h000000FFFFFFFFFFFFFC18000000003FFF00FFFFFC1EFFFFFF000000FFFFFFFF;
defparam sp_inst_9.INIT_RAM_1D = 256'hFFFFFC1FFFFFFF000000FFFFFFFFFFFFFE08000100003FFF017FFFFE1EFFFFFF;
defparam sp_inst_9.INIT_RAM_1E = 256'h000033001FFFFFFFFFFC0EFFFFFF800000FFFFFFFFFFFFFF040001C0001FFF83;
defparam sp_inst_9.INIT_RAM_1F = 256'hFFFFFFFFFFFF8204000FC00FFFFFFFFFF01FFFF7FF800000FFFFFFFFFFFFFF84;
defparam sp_inst_9.INIT_RAM_20 = 256'hFFE7FF800000FFFFFFFFFFFFFFC1003FFFE00FFFFFC1FFE01FFFE7FF800000FF;
defparam sp_inst_9.INIT_RAM_21 = 256'h87FFFFC000001FFFFFFF800000FFFFFFFFFFFFFFE0007FFFF107FFFFC03F001F;
defparam sp_inst_9.INIT_RAM_22 = 256'hFFFFF8007FFFFF47FFFFE000001FFFFFFF800000FFFFFFFFFFFFFFF0007FFFF9;
defparam sp_inst_9.INIT_RAM_23 = 256'h0000FFFFFFFFFFFFFFFC01FFFFFF43FFFFE000000FFFFFFF800000FFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_24 = 256'h00000FFFFFFF800000FFFFFFFFFFFFFFFC01FFFFFF83FFFFE000000FFFFFFF80;
defparam sp_inst_9.INIT_RAM_25 = 256'hFFFFFFC1FFFFF000000FFFFFFF800000FFFFFFFFFFFFFFFE00FFFFFF81FFFFE0;
defparam sp_inst_9.INIT_RAM_26 = 256'hFFFFFFFFFFFF807FFFFFE0FFFFF000000FFFFFFF800000FFFFFFFFFFFFFFFF00;
defparam sp_inst_9.INIT_RAM_27 = 256'hFFFFE00000FFFFFFFFFFFFFFFFC03FFFFFE0FFFFF000000FFFFFFFC00000FFFF;
defparam sp_inst_9.INIT_RAM_28 = 256'h7FFFF8000007FFFFFFF00000FFFFFFFFFFFFFFFFC03FFFFF607FFFF8000007FF;
defparam sp_inst_9.INIT_RAM_29 = 256'hFFFFF00FFFFFF87FFFF8000007FFFFFFF00000FFFFFFFFFFFFFFFFE01FFFFFF0;
defparam sp_inst_9.INIT_RAM_2A = 256'h00FFFFFFFFFFFFFFFFF80FFFFFFC3FFFF800000FFFFFFFF00000FFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_2B = 256'h0007FFFFFFF00000FFFFFFFFFFFFFFFFF807FFFFFC3FFFF800000FFFFFFFF000;
defparam sp_inst_9.INIT_RAM_2C = 256'hFFFFFE1FFFF8000007FFFFFFF00000FFFFFFFFFFFFFFFFFE03FFFFFF1FFFF800;
defparam sp_inst_9.INIT_RAM_2D = 256'hFFFFFFFFFFFF01FFFFFF07FFFC000007FFFFFFF00000FFFFFFFFFFFFFFFFFE03;
defparam sp_inst_9.INIT_RAM_2E = 256'hFFF80000FFFFFFFFFFFFFFFFFF01FFFFFF83FFFC000007FFFFFFF00000FFFFFF;
defparam sp_inst_9.INIT_RAM_2F = 256'hFFFC000007FFFFFFF80000FFFFFFFFFFFFFFFFFFC0FFFFFF83FFFC000007FFFF;
defparam sp_inst_9.INIT_RAM_30 = 256'hFFFFE03FFFFFC3FFFC000007FFFFFFF80000FFFFFFFFFFFFFFFFFFC07FFFFFC3;
defparam sp_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFEFE03FFFFFC3FFFC000007FFFFFFF80000FFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_32 = 256'h07FFFFFFF80000FFFFFFFFFFFFFFFFFFF01FEFFFE3F7FE000007FFFFFFF80000;
defparam sp_inst_9.INIT_RAM_33 = 256'hFFFFE183FF000007FFFFFFF80000FFFFFFFFFFFFFFFFFFF81FDFFFE1E7FE0000;
defparam sp_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFE0FFFFFF003FF000003FFFFFFF80000FFFFFFFFFFFFFFFFFFFC0F;
defparam sp_inst_9.INIT_RAM_35 = 256'hF80000FFFFFFFFFFFFFFFFFFFF07FFFFF803FF000003FFFFFFF80000FFFFFFFF;
defparam sp_inst_9.INIT_RAM_36 = 256'hFE000003FFFFFFF00000FFFFFFFFFFFFFFFFFFFF83FFFFF00FFF000003FFFFFF;
defparam sp_inst_9.INIT_RAM_37 = 256'hFFFFC1FFFFC000FE000003FFFFFFE00000FFFFFFFFFFFFFFFFFFFF83FFFFE005;
defparam sp_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFE07FFF0080FE000003FFFFFFC00000FFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_39 = 256'hFFFFFFE00000FFFFFFFFFFFFFFFFFFFFE01FFC008CFF000003FFFFFFC00000FF;
defparam sp_inst_9.INIT_RAM_3A = 256'hE0001FFF000003FFFFFFE00000FFFFFFFFFFFFFFFFFFFFE003F8001FFF000003;
defparam sp_inst_9.INIT_RAM_3B = 256'hFFFFFFFFFFF00000311FFF800003FFFFFF800000FFFFFFFFFFFFFFFFFFFFE000;
defparam sp_inst_9.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFFFFFFFFF00000039FFF800001FFFFFF800000FFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_3D = 256'h8000007FFFFFF04E3EFFF7FFFFFFFFFFFFFFFFFC000007FFFF800000FFFFFFF0;
defparam sp_inst_9.INIT_RAM_3E = 256'hFFFF800073FFFF0000007FFFFFFE8606FFFFFFFFFFFFFFFFFFFFFF000603EFFF;
defparam sp_inst_9.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFC000F7FFFF000001F3FFFFFFB000FFFFFFFFFFFFFFBFFF;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[30:0],sp_inst_10_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b00;
defparam sp_inst_10.BIT_WIDTH = 1;
defparam sp_inst_10.BLK_SEL = 3'b000;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'hF0E000033F0FFF740176678992C1903D9D19FC31C0FF0FB31800C000F01FE0FF;
defparam sp_inst_10.INIT_RAM_01 = 256'hF02487C130DFF7F3FE00077DFFFFC1CE7DE5F4E0C1B916CC27F80A42BF00A36C;
defparam sp_inst_10.INIT_RAM_02 = 256'hE3F161DFE6154043268C2313DF13FF3F8103F003FF7EFA1F08C91941650D943A;
defparam sp_inst_10.INIT_RAM_03 = 256'hE1C63FF5BC909AED8F21DB5AC86503D4E0F374A013F8038700E0E7FF186B0F98;
defparam sp_inst_10.INIT_RAM_04 = 256'h5B9C1790300CE0E3061C79721E5003BD2131560B4B06983F90579817C7F18FC0;
defparam sp_inst_10.INIT_RAM_05 = 256'hD02B258DCFDF9D537617AF191CF0E18C000B9472B66BB7A1BDF2377F040BC292;
defparam sp_inst_10.INIT_RAM_06 = 256'hFFB7CCE10B58D9E61A8BF7C14BD8FCF8E1AF429D78F817A9C752864EA430A0EB;
defparam sp_inst_10.INIT_RAM_07 = 256'hE0B300FC03D5C0FF79CA59CF58D8FBC8DC76219424EDCC505F434400FC9AA9C0;
defparam sp_inst_10.INIT_RAM_08 = 256'hB95422809942366D2C1F001C95FC030819A96A50E0B698CF35419DA5C5C25FB9;
defparam sp_inst_10.INIT_RAM_09 = 256'h2411ECE19CDB7897B7C8D83BEE7601F61F00AF3E7C0324DDAAEA50E4A8761D32;
defparam sp_inst_10.INIT_RAM_0A = 256'h7FACD900ABC01A6113077ED0780CEB4B80A70E20F8075A39F0D02A990101CF21;
defparam sp_inst_10.INIT_RAM_0B = 256'h501B481469900E116BE000878F30EA2F10340CACAC54D46B9B6718F8196A301C;
defparam sp_inst_10.INIT_RAM_0C = 256'hF71166AA88B507AF5F750D252C39794DA0019F6C7DC716A8C23B8DA854C7BCFA;
defparam sp_inst_10.INIT_RAM_0D = 256'hE9EE2B60182B4C3795A0A9FF8436DCD816CE2AC525878667C719827BDE7D2E46;
defparam sp_inst_10.INIT_RAM_0E = 256'hA8893AF9A02011AB4A060183D05060514237EBD5B0E1F17D3E56319AC9C9205C;
defparam sp_inst_10.INIT_RAM_0F = 256'h395E0E68EE620553344DCF9711964CE4C7500E2461D51D5EFF32F76B1E8CE5C4;
defparam sp_inst_10.INIT_RAM_10 = 256'hE9F54F039993175DD343B78E58FDAFA24FA928CB2BE1DCE4215B09A7CA463733;
defparam sp_inst_10.INIT_RAM_11 = 256'h7DA12DCD81F0A3C7AADF41502D12ED62FDC88435FA5CF6D9201C64AA3D9DC7CA;
defparam sp_inst_10.INIT_RAM_12 = 256'h17B806189B7B8951251D9F014594904E3F635CDE32EBAE7CDD5BE8D9DCA1F7DD;
defparam sp_inst_10.INIT_RAM_13 = 256'h2F37D87D061AD1E24006D0390AA240FFCF7CC0EB177C8E8600CF16000AD2D797;
defparam sp_inst_10.INIT_RAM_14 = 256'h80996D276780003DE234FFE2FF1FF341F897B0E81BB5E0C541CFF40A55248000;
defparam sp_inst_10.INIT_RAM_15 = 256'h06F44D4295B07B4F24A81CE2000E11EF358732C0D1AD4E07D43B52226F67285B;
defparam sp_inst_10.INIT_RAM_16 = 256'h78F7DAC2AFE0128490712311602F2024D04946001FCC6672936CE0E64869F024;
defparam sp_inst_10.INIT_RAM_17 = 256'h168028E4A32A968F10CD79561FE3F6EE6357EE08E08109B0C24280137557EFD1;
defparam sp_inst_10.INIT_RAM_18 = 256'h66796C001F857291C073F61C37CF990F86FBB38FFC4D5045EA1542AC0F6749A4;
defparam sp_inst_10.INIT_RAM_19 = 256'hAFA723678603B0FDE92484662285630C3A06282AF3DFA4EF5599039CDE1A05A0;
defparam sp_inst_10.INIT_RAM_1A = 256'h7A1D86016BE6FF4988B21FDBCAC0D7EF4A2B7AA461B08C3DCAE3D80E305B9FE5;
defparam sp_inst_10.INIT_RAM_1B = 256'h6378B4DB000EB75D40F6C60EF4CE7FDA45805A0A5C94143C352C5C496F802D5C;
defparam sp_inst_10.INIT_RAM_1C = 256'hFAAC944EF70A461174F0EE801E1CB273BBC52FBCFAC888DF83FEC74F01E80195;
defparam sp_inst_10.INIT_RAM_1D = 256'h066E484C4900453A7E642316F81731896557E0013C13EABECC5B33C839491CCA;
defparam sp_inst_10.INIT_RAM_1E = 256'h721D705AB69EF8DB302E909941B17A8607A92F6C6D845F3DED9A3EEB7A9B1697;
defparam sp_inst_10.INIT_RAM_1F = 256'hA2EDB272CF168D5DD7579CFF274632FA1801ED2EAE5FFF11152E59EB87C17B2F;
defparam sp_inst_10.INIT_RAM_20 = 256'hCC5410DFFF09E92DE8B4848F8887CD24397D0FB93CDE534B2DBB49B0DFFF0907;
defparam sp_inst_10.INIT_RAM_21 = 256'h34FF2E1908CA723FC982BFFF812161C357FD41781D830BB0C9CC66D0898F24DE;
defparam sp_inst_10.INIT_RAM_22 = 256'hC147150CE9550F777FB4E8F0043720DF20B5FFC1829AC40108FF07F89FC8BA85;
defparam sp_inst_10.INIT_RAM_23 = 256'hFFE9415732C5A097F7BE69F101FAE4F0170E00E8B0A129BCD5FFC95E4E0CADC0;
defparam sp_inst_10.INIT_RAM_24 = 256'h10342E5F3EDF35FFF98013282141688BE6AF7D58438C7FB71DB3384C4EDE4475;
defparam sp_inst_10.INIT_RAM_25 = 256'h67B0B3BAE0FCA4403F0D063FD4E2FFFB603DE932B79BC5759F6F7A36460065D0;
defparam sp_inst_10.INIT_RAM_26 = 256'h1C8E6BE93245751EC04489E3FCCE402444F355B0D3FFF9917C99862C0E4DEF11;
defparam sp_inst_10.INIT_RAM_27 = 256'h0D4762FFF08FE1FFE2C232A32EED604842ABBCE021B03225735C6F9FFFF9374C;
defparam sp_inst_10.INIT_RAM_28 = 256'h7516C54C087503016B7BFFF000231ED35B6CEB8C074A8B3CA545557DC81C6F70;
defparam sp_inst_10.INIT_RAM_29 = 256'hB91FC004F42E9779D8D8A41C1C003D1265FF702EC6006F0CB059D3A1A00FC847;
defparam sp_inst_10.INIT_RAM_2A = 256'h604FF81FD1E5BD7FFA102D840C2D531C5C181C5480993E43FF60557A1FF90481;
defparam sp_inst_10.INIT_RAM_2B = 256'h1E9A80D59DF483F03FE2FC44FA767B3C32585560D8FB38363019DA3F9F219BFF;
defparam sp_inst_10.INIT_RAM_2C = 256'h3F24BB76FE1FE8129501DFD6830F786D03CE90DCBBC697D33C1E0F95036068A4;
defparam sp_inst_10.INIT_RAM_2D = 256'hCE3A645FC27C78FB0E2BCC5A15880C8A4F5CDC983F183A367FA68796607CF17C;
defparam sp_inst_10.INIT_RAM_2E = 256'hE6F207180FE3C1817A727EE56DCDBC00907C422A4818045187CD821818263F16;
defparam sp_inst_10.INIT_RAM_2F = 256'h86AE981E1C9EB3D60B80F836AB6BB4FA1DDE83CB218A327E1D14ACB818046A17;
defparam sp_inst_10.INIT_RAM_30 = 256'hF36F37AF6C6A97A4A8180E2C7341586830F82C714546D1DACD7E8CF4CE424884;
defparam sp_inst_10.INIT_RAM_31 = 256'hFC0046B52C5988DF155492098539E926080C24B75BDABEEC7812FFECF25D90FB;
defparam sp_inst_10.INIT_RAM_32 = 256'h38CBF559EEFCE06FBE1C5EF75493EEFFB601974EE587A30E0A25CA155E62720E;
defparam sp_inst_10.INIT_RAM_33 = 256'hF7845B564AE00E7D0EE69AE13864C976FEAD5E18D6EC4E9479028EAE5075BC0A;
defparam sp_inst_10.INIT_RAM_34 = 256'hE8862F2BE4FFB58651DF933A4005FCFC5FFB981B521D884DA43FA4460A5C7812;
defparam sp_inst_10.INIT_RAM_35 = 256'h834582A019D7A4C8661AE247B64563D9810CCEEC0FD500680F50CA27A0C02104;
defparam sp_inst_10.INIT_RAM_36 = 256'h9EC40059F884BA2C8DDE300C68F0F88CE84BF9EAD0DC8066A76D620746FF8BC6;
defparam sp_inst_10.INIT_RAM_37 = 256'hFD6444BD6F085F2CCC06173153D908F1B6F4A234B2D7B13402FCD6ECFAF840DB;
defparam sp_inst_10.INIT_RAM_38 = 256'h2DA32688D3D8A7C8245338A68C5EBA7203DC1C75A88B0541C11BC0AA0DB2B923;
defparam sp_inst_10.INIT_RAM_39 = 256'hECBD03948F970BF5CE9CBEDA7C874F5C7A71F616BF787006E0E3B58317627C89;
defparam sp_inst_10.INIT_RAM_3A = 256'h4DF1A25D9806850D7282F8987C035F686E9B254ADE784EFC02B4824DAA980292;
defparam sp_inst_10.INIT_RAM_3B = 256'hED9CD0A6C680C6A144C5BBC8051013658E9A24F21E9B0F0F711BEA7DC4A3424A;
defparam sp_inst_10.INIT_RAM_3C = 256'hFA31E425CF57A4D8712908FFC60DFE02AB64AB0131AA14874EE56CBF5AD0CACB;
defparam sp_inst_10.INIT_RAM_3D = 256'h77FD8EE692B4A6D8251E717EDE8065784302AD948BDA8BCE1E4501E1F31F7431;
defparam sp_inst_10.INIT_RAM_3E = 256'h6CC03A939B8D0A9AA4AFCDEEAA2D920F1798334A144487BC57CC0A8D4F0D7046;
defparam sp_inst_10.INIT_RAM_3F = 256'hFB27B28ED2C097C00BF4AA7BE27CDDA320770F9CDF867BFEE3154AF8D92C37B6;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[30:0],sp_inst_11_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b00;
defparam sp_inst_11.BIT_WIDTH = 1;
defparam sp_inst_11.BLK_SEL = 3'b000;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'hFFFFFFFCC0F0FF3D000278FEA100D2B26CC2FFDE7FFF20241FFFFFFF0FE0FFFF;
defparam sp_inst_11.INIT_RAM_01 = 256'hFFC9FF00EF1407FFFFFFF88000FF890E034C8E5900B81E33E4FFEC7FBF2F340F;
defparam sp_inst_11.INIT_RAM_02 = 256'hC859803770ADBDFC34FCDF0C14E3FF3FFEFC0000FFCD9400D213D980BB93FDFD;
defparam sp_inst_11.INIT_RAM_03 = 256'h01C1FFEE3410795CB1C03B30F098FC98E0F08837E3F803F8FF00E0FF01AE0072;
defparam sp_inst_11.INIT_RAM_04 = 256'h9C1BE78FC0F01F0301FF76541E3F5543C0101FC502F820000F87EFE7C001F03F;
defparam sp_inst_11.INIT_RAM_05 = 256'hE44BBE71803F019B79E79FE1E00F0183FFB056FE88422EC0118B4B7EF8403FF3;
defparam sp_inst_11.INIT_RAM_06 = 256'h003FD865DB603607BD070500C7E5B7FF019F7CE100006077004FBE4048C1C020;
defparam sp_inst_11.INIT_RAM_07 = 256'hFF3C00009141C000E5DC18E3603706E44D04C04C3EB7CFE03F7C7800000680C0;
defparam sp_inst_11.INIT_RAM_08 = 256'h20CC3CD781C0F9F3CF1F002D2AFC0063FA2F0360175B0D9806604C3E97C3E07F;
defparam sp_inst_11.INIT_RAM_09 = 256'hE7A01B016A5600D86FF30F03A079FFC71F0099F8FC00293BCDD360134753B403;
defparam sp_inst_11.INIT_RAM_0A = 256'h910738008C628C9F40F08B6C9730CC27F4B70F5FBFFF633FF02300780019E42E;
defparam sp_inst_11.INIT_RAM_0B = 256'h6047BFF0721FFEF88F200038D14C0690F7C770079067338B9378473FF9733FFC;
defparam sp_inst_11.INIT_RAM_0C = 256'h0921403378E3F7CF803701C6339308D76001F85184A379E702B95A9067303793;
defparam sp_inst_11.INIT_RAM_0D = 256'h0EE50D865A1B8F28266031FF23C71F78B600CC7DCCFD96E0C7E1099BC1CF1F87;
defparam sp_inst_11.INIT_RAM_0E = 256'h30E269F60AE01E33FAA92F38309F0A64A2380C6DC3FEAE9CC09850FFEBD4E05F;
defparam sp_inst_11.INIT_RAM_0F = 256'hD2C1AB701FDEF963E3D94C6FF0186FFD5CF30DE0BE0B263EFF240FB2E05FDCF8;
defparam sp_inst_11.INIT_RAM_10 = 256'h42067084FD67F369BF55D8013F06CFE6A7A03838333F1D5690D201380A5B3FF0;
defparam sp_inst_11.INIT_RAM_11 = 256'h0E9E36DB00ED762ECCE080042BF6F62256130206FC9FF48BB0781CCCC4E35B36;
defparam sp_inst_11.INIT_RAM_12 = 256'hAE8A071F99D3C81699E954FE5668826BC081D49CF6F36057E985F2211FE52CC0;
defparam sp_inst_11.INIT_RAM_13 = 256'hA777DF7E07A1E5BB35F8E039E3B2E4FF982BFFF30DE77500000E5DFF0CCC981B;
defparam sp_inst_11.INIT_RAM_14 = 256'hFF9E652B220000456A07FF0ABD15B5CA00E7305CA8A2FF6BD7FFF83B96730000;
defparam sp_inst_11.INIT_RAM_15 = 256'h4BE835E119CAE77007F6273A000017AF06FFD4851AC63407E7412C75F078B537;
defparam sp_inst_11.INIT_RAM_16 = 256'h5625130160001CD59CCAB81A951F3F075A750600003E46040FBA150B7A11FFC7;
defparam sp_inst_11.INIT_RAM_17 = 256'hAD0018161D338B2225F68031E00327442328F4EA20FF0E399F3B000FE0BA0BCE;
defparam sp_inst_11.INIT_RAM_18 = 256'h87942000E033403A0010F132C735C52A7B0070F0006C8A03F0E65660FFF85340;
defparam sp_inst_11.INIT_RAM_19 = 256'h1460C085FC074001E76388991C2E000016028AE60644E5AEC1C500631AF80340;
defparam sp_inst_11.INIT_RAM_1A = 256'h8536FE5777B22B4BA7DEE26401E0C8E7390C829F0562001409F6CAF6979E76E0;
defparam sp_inst_11.INIT_RAM_1B = 256'hB428426B001A277FD7FE569B9B97B368537DE5FE834F0C0506C8CC3121401493;
defparam sp_inst_11.INIT_RAM_1C = 256'hC58C66E0F006C4582FBEC8600A28122B76545D9F7910F74D7DC5C36F51180486;
defparam sp_inst_11.INIT_RAM_1D = 256'hD99FFD80B68D3E05FFF85C0EF8FA40A12C50901428552474520D7F6FC1B68D3C;
defparam sp_inst_11.INIT_RAM_1E = 256'hD834FF09CC035A19FFD0D0F6CC8E857FE0AE1B700A04C08A864C15F3CFFAFB5D;
defparam sp_inst_11.INIT_RAM_1F = 256'hF90A2403FF31A9647070DAFFE4817F37D9774B6A808000E0461591F6073FAF02;
defparam sp_inst_11.INIT_RAM_20 = 256'h3C63480000F0A2F40AD8877F582E75B3674DBF81C3C301E8686854700000F0A5;
defparam sp_inst_11.INIT_RAM_21 = 256'hF800CF66CE0CD9C008564000785D740967FE3C2843B98880785C18EFF9AE28CA;
defparam sp_inst_11.INIT_RAM_22 = 256'h2B106EDE96B6DB5E00D87171B097C01F6B42003823F61201FF0AAF86DFB70C3E;
defparam sp_inst_11.INIT_RAM_23 = 256'h00109E676B963F5F505E4D46F12008F0DBA8B04018C0C87462003080815A9EFF;
defparam sp_inst_11.INIT_RAM_24 = 256'h8016629FC148A20000DFA46FB25E38581B026AA8675F003B4B40005071E1CCE2;
defparam sp_inst_11.INIT_RAM_25 = 256'h0DCFDFEF0000FA80123B0700334100009FA9574C98B8ACA8593848BBA3008637;
defparam sp_inst_11.INIT_RAM_26 = 256'hE3FC9AA6466E97A3FF685F83004680162503636FF800002FAAE7F4D1586D644E;
defparam sp_inst_11.INIT_RAM_27 = 256'h0320AC00005F22008CCA9380CE4B89CF94E4900094C00C778365DF9800005062;
defparam sp_inst_11.INIT_RAM_28 = 256'h284224080072FC00E7200000009B006CB0209B4330EB8CD792F79C9D70006180;
defparam sp_inst_11.INIT_RAM_29 = 256'hF418DAC7FDCE627E4A2150007400C309C20000B05700DF5B6FAD29AF2B0AEF3C;
defparam sp_inst_11.INIT_RAM_2A = 256'h00AA0000145EB3B6BE4140720C0E5E8EA9700E1BFFE40A7C0000A6430007A3AF;
defparam sp_inst_11.INIT_RAM_2B = 256'h0C1C001B88F8000096010389A101B07C7E242DE02C468AC2F00A1E3F1F143C00;
defparam sp_inst_11.INIT_RAM_2C = 256'h2707C76A5D06E80C190010CDC00080180331A545002EED7B31060F1AC8511710;
defparam sp_inst_11.INIT_RAM_2D = 256'h9D7CA61F9BC2C1530F3DEF9AF8F00013C0983BC800E091C700B2BABACF344280;
defparam sp_inst_11.INIT_RAM_2E = 256'hFE0A00E000E1C4BD3CE49FC21215610363328615700017CE05C3E407E0432B01;
defparam sp_inst_11.INIT_RAM_2F = 256'h0191020017BB921905000003ADE27ABC699F8517876509D86A136B3C0017DCF5;
defparam sp_inst_11.INIT_RAM_30 = 256'hFF09AE3CCE1F62C3A702000739116FF6C000141BD6CD7D043ECF8A45A5E98D26;
defparam sp_inst_11.INIT_RAM_31 = 256'hFA1B752D5F8B455F262A90DAF1F0B72F02000F7EEB1376F000071BB60F7E55D4;
defparam sp_inst_11.INIT_RAM_32 = 256'h27CCF367FEFF1CE0DC4B2828E1477F3085EB208E4DD351FC043ECCF3618EFC00;
defparam sp_inst_11.INIT_RAM_33 = 256'hC50453C7F940072B0F01E6003FE6C46BBA7675D58541F10B3CB30E53C42EC004;
defparam sp_inst_11.INIT_RAM_34 = 256'h1905E087BCF693C880C9C178A00D36006007611CCC1D00D678016A6DFBC389F6;
defparam sp_inst_11.INIT_RAM_35 = 256'h8ED9F63F636A7B26BBBC467FF05AE600D362CCB00736FFB000D133EF3F3D14FB;
defparam sp_inst_11.INIT_RAM_36 = 256'h5FF80031FFD77C0AA1A53F19074726D0AD78F96C6C8F00084772BC0037FFD3C7;
defparam sp_inst_11.INIT_RAM_37 = 256'h0188AF5D90A4B3F2000039FE843DF2AEA2FDDA90067AE379F9FFF437DD004906;
defparam sp_inst_11.INIT_RAM_38 = 256'hF05CC20F12603D1763C1239148929780013EFF666CF15205F9F2050CE31C863A;
defparam sp_inst_11.INIT_RAM_39 = 256'hE13E0367DAB090AAF816291DD466382D3DEC2AE2C4DA00021E1CC67BE433E453;
defparam sp_inst_11.INIT_RAM_3A = 256'hF8A1E8BB800209FE738300046F0B2B9F6FC5C35CA5F814ED2F1A01BBD1C00603;
defparam sp_inst_11.INIT_RAM_3B = 256'h13301F2FE83DB186388059F0030A0C99730410D51393F12E43E004814FD07BB4;
defparam sp_inst_11.INIT_RAM_3C = 256'h417D596BFCBF24C57D0F3FE184C4F9FFD2704C001066188280AD282287FB710F;
defparam sp_inst_11.INIT_RAM_3D = 256'hD603CDB736AE164C80BF956433DC61D7DC7D5ACFA6B1136FC056002455280EA1;
defparam sp_inst_11.INIT_RAM_3E = 256'h4667C1A6EA9E3A103C5E40182829FC1EB04B3343B080E56B3E7E5683EB14CEFF;
defparam sp_inst_11.INIT_RAM_3F = 256'hB6657DF1192D4DFA60D2A44B2CAB7F3CD74A6701C4279339C0C063E010CB0400;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[30:0],sp_inst_12_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b00;
defparam sp_inst_12.BIT_WIDTH = 1;
defparam sp_inst_12.BLK_SEL = 3'b000;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFFFFFF03FFFEDF00AA0071C40868001F7F00E0381FFFFFFFFFFFFFFF;
defparam sp_inst_12.INIT_RAM_01 = 256'h000EFFFFE01807FFFFFFFFFFFFFF06F1FF23C06A0068E4044C000F7F40E0380F;
defparam sp_inst_12.INIT_RAM_02 = 256'hB06A000D00C0540038FCFF001803FF3FFFFFFFFFFFAC0FFFC9E06A0017620654;
defparam sp_inst_12.INIT_RAM_03 = 256'hFE3FFFE533EFF8C1AA000601E65400E0E0F0003803F803FFFFFF1FFF1591FFF6;
defparam sp_inst_12.INIT_RAM_04 = 256'h1FE0078000FFFFFCFFFF70D0E1FF31EA000FC622D600C0000007F007C001FFFF;
defparam sp_inst_12.INIT_RAM_05 = 256'h51C42A010000FE1C80078001FFFFFE7FFF800E017FC6CB000EA3B86A0080000C;
defparam sp_inst_12.INIT_RAM_06 = 256'h00703FFD18800FEF988906003FFE3800018080FEFFFFFFFF004681BFFB85001F;
defparam sp_inst_12.INIT_RAM_07 = 256'h003FFFFFF0D6C000543FE7FD800FF7E58707003C3F38300000807FFFFFFE8FC0;
defparam sp_inst_12.INIT_RAM_08 = 256'hC03C3F187E3F00000FE0FFE39BFC000906D0FC800FEFEE4707803C3F183C0000;
defparam sp_inst_12.INIT_RAM_09 = 256'h18C007FCFEA900E01FFC10FC60800007E0FF5F64FC002307F03C800FFBB34F03;
defparam sp_inst_12.INIT_RAM_0A = 256'h4567F8008F519000600FF16C6900F01FF8B8F0C0C00083C00FA464F800194330;
defparam sp_inst_12.INIT_RAM_0B = 256'h80C0400F83E0014260E0003F55C801200FF8A2BD80780FF39C80C0400683C003;
defparam sp_inst_12.INIT_RAM_0C = 256'h303DC03C073FF80F4048FE07C008F898E001FF8C5080A01FFC75BD80780FC79C;
defparam sp_inst_12.INIT_RAM_0D = 256'hF0E360809DFBF0083BE03E003FF81F38C9FF0F825C23D9E0C7FE0790C010FFF8;
defparam sp_inst_12.INIT_RAM_0E = 256'h3F1E70CC43E01FC3F9A2A0C3F0E0107AE23FF07DFCFF9F03FF1F8FC123C7E05F;
defparam sp_inst_12.INIT_RAM_0F = 256'h1C3FCC7FFFC1FE7C1CEBB830F01F8FFCB13191E0C00C39FEFF38003CFFC0C3FF;
defparam sp_inst_12.INIT_RAM_10 = 256'h35078000DEBFF08E7F661FFF00F8F01ECFD008F83C3F1C8ABBBC01C0039C7FF0;
defparam sp_inst_12.INIT_RAM_11 = 256'h597FC738FF1E9FED0F0002E797F107E267E3FEF800E00F0CE00DFCF0FC00256C;
defparam sp_inst_12.INIT_RAM_12 = 256'h3D8C07E06633A01A7E0E33FFD8DB878C0000A742F103E067F1FCFC01E01C1EE0;
defparam sp_inst_12.INIT_RAM_13 = 256'h3A9C208007C006390600FFC61CD8490010E7FFFC4185D80000F2A400F0C0E01C;
defparam sp_inst_12.INIT_RAM_14 = 256'hFF9F90421800000999F8000D3CE63333FF07CF801E6F0070CFFFFF80A6880000;
defparam sp_inst_12.INIT_RAM_15 = 256'h8E4036B5E1061F7F0748B2CC000020D8F80018FCE302F807F87F401A0980C30F;
defparam sp_inst_12.INIT_RAM_16 = 256'h64ECE3FF1FFFE0E42023F2E30CFF3F07A4B0A400001559F800330CF386FE0007;
defparam sp_inst_12.INIT_RAM_17 = 256'h360007F220C383CBEC07FF0FFFFC38781CF00719E0FF0FC6192000001409F3C0;
defparam sp_inst_12.INIT_RAM_18 = 256'h07F3E000FFFE4432000FF206070616E603FF0FFFFF8EFC000107B1E0FFFFED0A;
defparam sp_inst_12.INIT_RAM_19 = 256'hFC1FFFF980000001E0E070FFFF8E6B000E01361E0468229499C2FFFFE3840000;
defparam sp_inst_12.INIT_RAM_1A = 256'h48F20498E3E1B7B79FE1FC000700C0E0F8F0FD7F65DC000C08F9C604D852ECC1;
defparam sp_inst_12.INIT_RAM_1B = 256'hC718FEDC4006388832049987F7EC00D860FE0006E0C003FCF8F03C79AC800C1F;
defparam sp_inst_12.INIT_RAM_1C = 256'h0073F8DF0FFE389F1F48974006300519049B2F3FFBC0506CFE003F70CE07FC78;
defparam sp_inst_12.INIT_RAM_1D = 256'h5BFFFA20502CFFC000003FFEF8037F9E906B200C30761DF89E7CFFFD21502CFF;
defparam sp_inst_12.INIT_RAM_1E = 256'h9C0CFF9C020399D4FFFB30506C7FC000006FF8800CFBC0093B900CFC2A06039C;
defparam sp_inst_12.INIT_RAM_1F = 256'h17F3C7FC00F041863070ED00E700D9FFFA8927B67FC00000C7F3E1FBF8FFBE1B;
defparam sp_inst_12.INIT_RAM_20 = 256'h0380C7C000006313F31F7800C7EC86904078C07E003E3E5C9E18630FC0000066;
defparam sp_inst_12.INIT_RAM_21 = 256'h2400F00030F03D000831C00000C193F27800031837C258DF7A63FF0006907033;
defparam sp_inst_12.INIT_RAM_22 = 256'h18CF835050271805FF1F1B7E7875001F18C000009CF1E4FE0006601EE2502F3D;
defparam sp_inst_12.INIT_RAM_23 = 256'h0000BF874C48C030CFDE83D021C796F0E3A5C0307200080CC00000BF00937F00;
defparam sp_inst_12.INIT_RAM_24 = 256'h000810E00038800000BFC7B09360E7C7D8A898287FD0003C0080003280003CC0;
defparam sp_inst_12.INIT_RAM_25 = 256'hD2001F5E0000E8000C05F800F0C00000BFCE60202087638059B8683EEA0007C8;
defparam sp_inst_12.INIT_RAM_26 = 256'h00A0A6608E77BE90008F7F830050000801FC80E0A000009FCC00A8A3389AB7EC;
defparam sp_inst_12.INIT_RAM_27 = 256'hFF1FD80000C03400A0798CC00E5E0030181F10001E00001EFC83C0300000CF8B;
defparam sp_inst_12.INIT_RAM_28 = 256'hDF9E07700007FF001F24000000D300DFF71F2CC0FB2270E78FC81C1E800016FF;
defparam sp_inst_12.INIT_RAM_29 = 256'hD0BD27A6060E019F96037800040000F81C00003F67003FC71FD9A25DB2F30F03;
defparam sp_inst_12.INIT_RAM_2A = 256'h00330000133F6FD17CB3FC040C0DDFD2037800000003F99C0000388300009F9F;
defparam sp_inst_12.INIT_RAM_2B = 256'h0003FFE07B1C000024000004622FD6FE9F2009E00DBFD609F80401C0E0F3DC00;
defparam sp_inst_12.INIT_RAM_2C = 256'h3707FF886308100002FFE03C1C0000500300933917A1FFC2E5160F1EAF9F08F8;
defparam sp_inst_12.INIT_RAM_2D = 256'hBCFF827FEC3D0A630F3B1A19FE0000003FE007E400002007006E7C36DFF93FE0;
defparam sp_inst_12.INIT_RAM_2E = 256'hFE08000005F5C37CFF1DFFC03DA14100F7AFFEFE8000043FF9C00C0000813300;
defparam sp_inst_12.INIT_RAM_2F = 256'hFF86FC00047C8C1F0A00000A45E6FE7FEBFF513AFC41073520EF16C000043F09;
defparam sp_inst_12.INIT_RAM_30 = 256'hDFCE07C1DAEE64FFA6FC0014FDCE8FFB000009E9CDC83E5D5F5F0C98C1D8B183;
defparam sp_inst_12.INIT_RAM_31 = 256'hF2E92CC93F0783FFF80C6DCDB1673F26FC0014FB24E3FB00000AE9920BC09330;
defparam sp_inst_12.INIT_RAM_32 = 256'h1430F0800B0000E5E838F21FD170DF608333630E51F1CE00001430F0800B0000;
defparam sp_inst_12.INIT_RAM_33 = 256'h89047E053B80001CF00001F5C018C37179FA7331F3DEA00371F40E5ED11C0000;
defparam sp_inst_12.INIT_RAM_34 = 256'hB3061F3FC30157F000EF82FAC00209FF8000F5E03F1D05DDFDB4E36304600443;
defparam sp_inst_12.INIT_RAM_35 = 256'h8BC10E3FD754FDAA3C7F7E7FFFF20000E60CCEC00009FFC00025FC1F3FEB21FD;
defparam sp_inst_12.INIT_RAM_36 = 256'h6200000FFFE7FFF39EC33F44523AAAE06E780690A6000024077DC00009FFE3C7;
defparam sp_inst_12.INIT_RAM_37 = 256'h0180D41A00A0034200000FFFE7FE039F01FCB9277B763FFE07FFF7A8C0004030;
defparam sp_inst_12.INIT_RAM_38 = 256'hEEF8FE0F1668C31FE026260100842200000EFF87EF02CFA2FBF4F270E0227FC6;
defparam sp_inst_12.INIT_RAM_39 = 256'h1E3FFC07C3CFB7D7FFEDCF1BCCBDF80C8AC9E320F56580010EFF07FC07EC43C8;
defparam sp_inst_12.INIT_RAM_3A = 256'h7918670640010000737C00079F5BAFFF9A1700FFC3D7EA6D1D9084A0A680010D;
defparam sp_inst_12.INIT_RAM_3B = 256'h007A1FAFF9010820608CC6C000020001FC000737B3FFF8E56B00A5010FE9FA03;
defparam sp_inst_12.INIT_RAM_3C = 256'h3D01C1B5E7AF30C3E90FB7F7FB6200173E8330000BE1E0830096EF63F5E9D71B;
defparam sp_inst_12.INIT_RAM_3D = 256'h98003392D94026398180340A53E863F7C02BEE01D00039F0C018001C333000C1;
defparam sp_inst_12.INIT_RAM_3E = 256'h7DDA1841A01FBB1FC34039EFD3EE092A8FF47EE3D802D6E7F51222200C750C7F;
defparam sp_inst_12.INIT_RAM_3F = 256'h86E64002B87E4C0622D4445CBFA57EC04F8408013CE7683FE3472340E2A8CCDD;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[30:0],sp_inst_13_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b00;
defparam sp_inst_13.BIT_WIDTH = 1;
defparam sp_inst_13.BLK_SEL = 3'b000;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h00000000000000FFFFFE3FFF4C003007F027FFE07FFFE03FE000000000000000;
defparam sp_inst_13.INIT_RAM_01 = 256'hFFF0FFFFE01FF800000000000000FFFFFF1FFF8C001807F823FFF07FFFE03FF0;
defparam sp_inst_13.INIT_RAM_02 = 256'h7F8C000300FE33FFC0FCFF001FFC00C0000000000033FFFFC7FF8C000F03F833;
defparam sp_inst_13.INIT_RAM_03 = 256'h00000019CFFFF83E4C000100FF33FF00E0F0003FFC07FC0000000000E67FFFF1;
defparam sp_inst_13.INIT_RAM_04 = 256'h1FFFF87FFF00000000008F6FFFFF0E0C0000C60F31FF00000007FFF83FFE0000;
defparam sp_inst_13.INIT_RAM_05 = 256'h3157D9FE0000001FFFF87FFE00000000007FE9FFFFC10C0000630F99FF000000;
defparam sp_inst_13.INIT_RAM_06 = 256'hFF4FFFFD1A00001F93F8F80000003FFFFE7FFF0000000000FFBB7FFFF8060000;
defparam sp_inst_13.INIT_RAM_07 = 256'hFFC000000FD83FFF9BFFFFFE00000FE1FCF80003C03FFFFFFFFF80000001703F;
defparam sp_inst_13.INIT_RAM_08 = 256'h0003C01FFFFFFFFFF000001F6C03FFF2FEFFFF000007E9FCF80003C01FFFFFFF;
defparam sp_inst_13.INIT_RAM_09 = 256'hFF000003FDF8FF0000001FFFE0FFFFF800003FF703FFDDFFFFFF000007F1FCFC;
defparam sp_inst_13.INIT_RAM_0A = 256'hC60807FF709F9FFF800000ED78FF000000BFFFC0FFFFFC000067F707FFE67F3F;
defparam sp_inst_13.INIT_RAM_0B = 256'hFFC07FFFFC0000C3F01FFFC026CFFFC00000623C7F8000039FFFC07FFFFC0000;
defparam sp_inst_13.INIT_RAM_0C = 256'h103C3FC0003FFFF0C07FFFF80007F8E01FFE0001C77FC00000313C7F8000079F;
defparam sp_inst_13.INIT_RAM_0D = 256'h00E0B97FE00400183E1FC0003FFFE0F8FFFFF0003C3FE01F380000F33FE00000;
defparam sp_inst_13.INIT_RAM_0E = 256'hC00101E8231FE003F84EDFFC0F00087E1DC0007DFF007FFFFFE00040CC381FA0;
defparam sp_inst_13.INIT_RAM_0F = 256'hE0000F80003FFF80020ED0100FE00FFC074F9E1F00043F0100C0003F003F3FFF;
defparam sp_inst_13.INIT_RAM_10 = 256'h07F800021F800FF00087E000FFFF000309201807C03F1C03A79FFE00061F000F;
defparam sp_inst_13.INIT_RAM_11 = 256'h1D0007F80000F917F0000107800FF81D87FC01FFFF00020FC0210300FC0001F2;
defparam sp_inst_13.INIT_RAM_12 = 256'hC38FF800000C707A000FF000207C7BF0000087C10FFC1F87FE03FFFE0003FF00;
defparam sp_inst_13.INIT_RAM_13 = 256'h63F3FFFFF80007C707FF0000004317001FE000001E39E0000043E3FFFF3F001F;
defparam sp_inst_13.INIT_RAM_14 = 256'h006007BC70000021F7FFFFF03C07CF03FFF800005CE9007FC000000F58F00000;
defparam sp_inst_13.INIT_RAM_15 = 256'hF180178601FE0080F803DC70000010F7FFFFE0FC03FE0007FF80802C0F00FF00;
defparam sp_inst_13.INIT_RAM_16 = 256'h871C03FF000000FBC01C7C03FC00C0F801C63800000C77FFFFC3FC03FE000007;
defparam sp_inst_13.INIT_RAM_17 = 256'h3800000E3BFC7C0C1C07FF0000003F80000007F81F00F000E23C00000C3FFC3F;
defparam sp_inst_13.INIT_RAM_18 = 256'h07F01FFF0000FBBC00000E1DF8F8181E03FF0000000F00000007F01F00000075;
defparam sp_inst_13.INIT_RAM_19 = 256'hFC00000100000001E01FFF000051AE0001FF3E01F8701E78C1C0000003000000;
defparam sp_inst_13.INIT_RAM_1A = 256'hCFF1F8E017C03FFF800000800000C0E007FF00008A9F0003F7FFC1F8E029F721;
defparam sp_inst_13.INIT_RAM_1B = 256'h0707050F8001C04FF1F8E06F0FF7FFC78000800100C00003FF00038E0F0003E0;
defparam sp_inst_13.INIT_RAM_1C = 256'h800000C00001FF1F0003278001C047F8F8E0FE7FFE3FCF8C00800080C00003FF;
defparam sp_inst_13.INIT_RAM_1D = 256'hFCFFFE1FCFCC00800000000107FC7F800193C003C037FC00E1DEFFFC1ECFCC00;
defparam sp_inst_13.INIT_RAM_1E = 256'hE0030009FE03E7F9FFF80FCF8C008000001007FFF0FFC009CBE003001BFE03E3;
defparam sp_inst_13.INIT_RAM_1F = 256'h0FFC07FFFFF075F80F8F04FFE7FFC0FFEC1EE03E00800000380FFE03FFFFBE63;
defparam sp_inst_13.INIT_RAM_20 = 256'hFFFFC08000001C0FFC1FFFFFC032F8707F84FFFFFFFEFF901FF87F0080000018;
defparam sp_inst_13.INIT_RAM_21 = 256'h3C00FFFFFF0011FFF7F08000003E0FFC7FFFFF07D9FCC71F867FFFFFFF804013;
defparam sp_inst_13.INIT_RAM_22 = 256'hF83FF4DFCFC7E71C001FE7800019FFE0F88000007F0FF8FFFFFE1FE9FCCFCFC3;
defparam sp_inst_13.INIT_RAM_23 = 256'h00007FF88FC0FFF03FE54FCFC1FF9D0F03B300001CFFF7FC8000007FFFE3FFFF;
defparam sp_inst_13.INIT_RAM_24 = 256'h00001CFFFFF8C000007FF83F8C7FE03FE36E07C87FDDFFC01000001CFFFFFC80;
defparam sp_inst_13.INIT_RAM_25 = 256'h60001F7EFFFF00000011FFFFF08000007FF07F1F3F801FF1BFC7883EEFFFF810;
defparam sp_inst_13.INIT_RAM_26 = 256'hFF9F3E1F0187CFE0000F7F7CFFA8000011FFFFE0C000007FF0FF9F3F0707C79F;
defparam sp_inst_13.INIT_RAM_27 = 256'hFF001000003FC7FF9F787F000E67B0001FFF6FFFE800000FFFFFC02000003FF3;
defparam sp_inst_13.INIT_RAM_28 = 256'hBFE1F080000FFF0000C80000FF1CFFC0F0FFCFC027D200F87FBFE3E800000FFF;
defparam sp_inst_13.INIT_RAM_29 = 256'hE77E09E607F1FFBFE1F480000C000007E80000C078FFFFC0FFEE9C13E203F0FF;
defparam sp_inst_13.INIT_RAM_2A = 256'h00C3FFFFEF001FE7FF04FC07F3F3FFE1F4800008000007E80000C0FCFFFF807F;
defparam sp_inst_13.INIT_RAM_2B = 256'h0008000007E80000C7FFFFFC1C1FE6FF04BC0E1FF3DFE1F400000800000FE800;
defparam sp_inst_13.INIT_RAM_2C = 256'h38F800E780F4000008000003E800009FFCFF70FE0FDFFE3E7D19F0E1FFE0F400;
defparam sp_inst_13.INIT_RAM_2D = 256'h83FF3E3FF0FEAE7CF0C7F818040000080000000800003FF8FFE1FF313FFEFD2C;
defparam sp_inst_13.INIT_RAM_2E = 256'hFE0C0000FC063F03FFA3BF80FED77EFFF0DFFE0400000C0001C0080000FF3CFF;
defparam sp_inst_13.INIT_RAM_2F = 256'hFF8400000C00801F0C0000F9F61E01FFB7BF8EFCCF7EFF0E5FFF0400000C0001;
defparam sp_inst_13.INIT_RAM_30 = 256'h3F8FF3FE39F1BCFFA400000C01C00FFC0000FBF23C30FF9C3FBFF0E5FE387E3F;
defparam sp_inst_13.INIT_RAM_31 = 256'h09F2E3F10000003FBFF2FE3BCEBC3F2400000C03E003FC0000F9F271F33F100F;
defparam sp_inst_13.INIT_RAM_32 = 256'h0C00F0000C00001C0F07FCFFCE703FBF797C17F19C1BC200000C00F0000C0000;
defparam sp_inst_13.INIT_RAM_33 = 256'h5EFB9E41050000040000000600003F7F07FC8F0EF03F3FFC5E1FF19E05010000;
defparam sp_inst_13.INIT_RAM_34 = 256'hC8F8003FFFFE44BFFF0F0204000004000000060000E2FC23FECC1C60007FFEF4;
defparam sp_inst_13.INIT_RAM_35 = 256'h8C3E01C0309DFED9C0007E7FFF3AFFFF040530000004000000060000C018C3FE;
defparam sp_inst_13.INIT_RAM_36 = 256'h830000040007FFFC7F00C0C39EFCD900107800008FFFFFC804810000040003C7;
defparam sp_inst_13.INIT_RAM_37 = 256'hFE7F2FE7FF0005830000040007FFFC7FC00387C7038E3F000000085F3FFF900A;
defparam sp_inst_13.INIT_RAM_38 = 256'h1FFD01F0EE6700E01FDF59FE804EC30000050007EFFC3FC0070FFBFF1F3E0001;
defparam sp_inst_13.INIT_RAM_39 = 256'h003FFFF83C00700FFD03F0E7C33C07F3D7261E005B810000050007FFF81F8038;
defparam sp_inst_13.INIT_RAM_3A = 256'h1030B0008000040073FFFFF800C427FD0618FFC0FFCFF1D3846400FCC0000004;
defparam sp_inst_13.INIT_RAM_3B = 256'hFF03E07FF0E2C0401AE0C08000060001FFFFF8088CF7FD1C8CFF99FEDFF0C581;
defparam sp_inst_13.INIT_RAM_3C = 256'hFEFE3E3C0860C73F0EF06FF838C0003C6200400007E00083FF78101CF3F230EC;
defparam sp_inst_13.INIT_RAM_3D = 256'hE0000071E00039F9817FDBF1CC0F9F183FE7F1FA60000250C0600003F0C000FE;
defparam sp_inst_13.INIT_RAM_3E = 256'h7C3C70090CBF3BE0003FFBF003EFF93B7FE801DC1FFE181FF3E1FCF0003E077F;
defparam sp_inst_13.INIT_RAM_3F = 256'h86187FFE27DF93FE1CE8032B9F2180003FFDF001FCE79C1FF4C71C7FFE37231C;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[30:0],sp_inst_14_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b00;
defparam sp_inst_14.BIT_WIDTH = 1;
defparam sp_inst_14.BLK_SEL = 3'b000;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h00000000000000000001FFFFF0000FF8001FFFFF80001FC00000000000000000;
defparam sp_inst_14.INIT_RAM_01 = 256'hFFFF00001FE00000000000000000000000FFFFF00007F8001FFFFF80001FC000;
defparam sp_inst_14.INIT_RAM_02 = 256'hFFF00000FF000FFFFF0300FFE00000000000000000C000003FFFF00000FC000F;
defparam sp_inst_14.INIT_RAM_03 = 256'h000000FE000007FFF00000FF000FFFFF1F0FFFC00000000000000000F800000F;
defparam sp_inst_14.INIT_RAM_04 = 256'hE0000000000000000000FF800000FFF0000039F00FFFFFFFFFF8000000000000;
defparam sp_inst_14.INIT_RAM_05 = 256'h0EB807FFFFFFFFE0000000000000000000FFF000003FF000001CF007FFFFFFFF;
defparam sp_inst_14.INIT_RAM_06 = 256'hFF800002E40000006C07FFFFFFFFC0000000000000000000FFFC000007F80000;
defparam sp_inst_14.INIT_RAM_07 = 256'h000000000020FFFFE00000000000001E03FFFFFFFFC0000000000000000000FF;
defparam sp_inst_14.INIT_RAM_08 = 256'hFFFFFFE00000000000000000F0FFFFFC0100000000001603FFFFFFFFE0000000;
defparam sp_inst_14.INIT_RAM_09 = 256'h000000000307FFFFFFFFE0001F000000000000F8FFFFFE0000000000000E03FF;
defparam sp_inst_14.INIT_RAM_0A = 256'h38F0FFFFFFE060000000001387FFFFFFFF40003F000000000018F8FFFFFF80C0;
defparam sp_inst_14.INIT_RAM_0B = 256'h003F80000000003C00FFFFFFF830000000001DC3FFFFFFFC60003F8000000000;
defparam sp_inst_14.INIT_RAM_0C = 256'h0FC3FFFFFFC000003F80000000000700FFFFFFFE38000000000EC3FFFFFFF860;
defparam sp_inst_14.INIT_RAM_0D = 256'hFF1FC60000000007C1FFFFFFC00000070000000003C000FFFFFFFF0C00000000;
defparam sp_inst_14.INIT_RAM_0E = 256'h0000FFF01CFFFFFC07F1000000000781FFFFFF82000000000000003FF000FFFF;
defparam sp_inst_14.INIT_RAM_0F = 256'hFFFFF0000000000001F1E00FFFFFF003F88060000003C0FFFFFFFFC000000000;
defparam sp_inst_14.INIT_RAM_10 = 256'hF8000001E07FFFFFFFF8000000000001F0C007FFFFC0E3FC4060000001E0FFFF;
defparam sp_inst_14.INIT_RAM_11 = 256'h3EFFF807FFFF00F8000000F87FFFFFFFF8000000000001F0001EFFFF03FFFE01;
defparam sp_inst_14.INIT_RAM_12 = 256'h007000000000003DFFF00FFFFF80FC000000783FFFFFFFF80000000000000000;
defparam sp_inst_14.INIT_RAM_13 = 256'h1C0FFFFFFFFFF800F8000000003C38FFE01FFFFFE07E0000003C1FFFFFFFFFE0;
defparam sp_inst_14.INIT_RAM_14 = 256'hFFFFF81F8000001E0FFFFFFFC3F800FC000000003F10FF803FFFFFF03F000000;
defparam sp_inst_14.INIT_RAM_15 = 256'h00000878FE01FFFFFFFC0F8000000F0FFFFFFF03FC01FFF80000001FF0FF00FF;
defparam sp_inst_14.INIT_RAM_16 = 256'hF803FC00FFFFFF00000000FC03FFFFFFFE0FC00000038FFFFFFC03FC01FFFFF8;
defparam sp_inst_14.INIT_RAM_17 = 256'hC0000001C7FFFFF003F800FFFFFFC0000000F807FFFFFFFF07C0000003C7FFFF;
defparam sp_inst_14.INIT_RAM_18 = 256'hF80FFFFFFFFF81C0000001E3FFFFE001FC00FFFFFFF0000000F80FFFFFFFFF83;
defparam sp_inst_14.INIT_RAM_19 = 256'h03FFFFFE000000FE1FFFFFFFFFE0D0000000C1FFFF8001FF3E3FFFFFFC000000;
defparam sp_inst_14.INIT_RAM_1A = 256'h300FFF000FFFC0007FFFFF0000003F1FFFFFFFFFF060000000003FFF0007F81E;
defparam sp_inst_14.INIT_RAM_1B = 256'hF8FFF830000000300FFF001FFFF8003FFFFF0000003FFFFFFFFFFFF070000000;
defparam sp_inst_14.INIT_RAM_1C = 256'h0000003FFFFFFFE0FFFC180000003807FF001FFFFC003FF3FF0000003FFFFFFF;
defparam sp_inst_14.INIT_RAM_1D = 256'h3FFFFC003FF3FF000000FFFFFFFF807FFE0C0000000803FF003FFFFE003FF3FF;
defparam sp_inst_14.INIT_RAM_1E = 256'h0000000601FC003FFFFC003FF3FF000000FFFFFFFF003FF6040000000401FC00;
defparam sp_inst_14.INIT_RAM_1F = 256'hFFFFF800000F82000000030018003FFFF0001FC1FF000000FFFFFFFC00004184;
defparam sp_inst_14.INIT_RAM_20 = 256'h00003F000000FFFFFFE000003FC1000F800300000001FFE0000780FF000000FF;
defparam sp_inst_14.INIT_RAM_21 = 256'hC3FF000000000E00000F000000FFFFFF800000FFE0003FE001800000007F800C;
defparam sp_inst_14.INIT_RAM_22 = 256'h07FFF8203FF800E3FFE00000000E000007000000FFFFFF000001FFF0003FF000;
defparam sp_inst_14.INIT_RAM_23 = 256'h0000FFFFF03F000FFFF8303FFE0063FFFC4000000F000003000000FFFFFC0000;
defparam sp_inst_14.INIT_RAM_24 = 256'h00000F000007000000FFFFC07F801FFFFC11FFF78023FFFFE000000F00000300;
defparam sp_inst_14.INIT_RAM_25 = 256'hFFFFE081FFFFF000000E00000F000000FFFF80FFC07FFFFE00FFF7C111FFFFE0;
defparam sp_inst_14.INIT_RAM_26 = 256'h007FC1FFFFF8007FFFF080FFFFF000000E00001F000000FFFF007FC0FFFFF800;
defparam sp_inst_14.INIT_RAM_27 = 256'h00FFE00000FFF8007F87FFFFF1807FFFE000FFFFF000000000003FC00000FFFC;
defparam sp_inst_14.INIT_RAM_28 = 256'h7FFFF800000000FFFFF00000FFE0003F0FFFF03FC03DFF00007FFFF000000000;
defparam sp_inst_14.INIT_RAM_29 = 256'hF8FFF019F800007FFFF8000003FFFFFFF00000FF8000003FFFF07FE01DFC0000;
defparam sp_inst_14.INIT_RAM_2A = 256'h00FC000000FFFFF8FFF803F800003FFFF8000007FFFFFFF00000FF0000007FFF;
defparam sp_inst_14.INIT_RAM_2B = 256'h0007FFFFFFF00000F8000003FFFFF9FFF843F000003FFFF8000007FFFFFFF000;
defparam sp_inst_14.INIT_RAM_2C = 256'hC000001FFFF8000007FFFFFFF00000E000000FFFFFFFFFFC02E000001FFFF800;
defparam sp_inst_14.INIT_RAM_2D = 256'h7FFFC1FFFFFF1180000007E7F8000007FFFFFFF00000C000001FFFCFFFFFFE13;
defparam sp_inst_14.INIT_RAM_2E = 256'h01F0000003F800FFFFC07FFFFF0880000F0001F8000003FFFE3FF0000000C000;
defparam sp_inst_14.INIT_RAM_2F = 256'h0078000003FF7FE0F0000007F801FFFFC07FFFFF008000FF8000F8000003FFFE;
defparam sp_inst_14.INIT_RAM_30 = 256'hFFF0000007FFC30058000003FE3FF000000007FC03FFFFE3FFFFFF020007FFC0;
defparam sp_inst_14.INIT_RAM_31 = 256'h07FC1FFEFFFFFFFFC0010007FFC3C0D8000003FC1FFC00000007FC0FFCFFEFFF;
defparam sp_inst_14.INIT_RAM_32 = 256'h03FF0FFFF0000003F0FFFF003F8FFFC000800FFFE3E43C000003FF0FFFF00000;
defparam sp_inst_14.INIT_RAM_33 = 256'h3FFFE182FE000003FFFFFFF800000080FFFF00FF0FFFC000800FFFE1E2FE0000;
defparam sp_inst_14.INIT_RAM_34 = 256'h07FFFFC00000287FFFF001FF000003FFFFFFF800000003FFFF03FF9FFF800008;
defparam sp_inst_14.INIT_RAM_35 = 256'h700000000FE3FF07FFFF81800005FFFFF803FF000003FFFFFFF800000007FFFF;
defparam sp_inst_14.INIT_RAM_36 = 256'hFC000003FFF800000000003FE1FF07FFFF87FFFF13FFFFF00FFE000003FFFC38;
defparam sp_inst_14.INIT_RAM_37 = 256'hFFFFC1FFFFC000FC000003FFF800000000007FF8FC01C0FFFFFFFF83FFFFE005;
defparam sp_inst_14.INIT_RAM_38 = 256'hFFFE0000019FFFFFFFE0FFFF0181FC000003FFF81000000000FFFC0000C1FFFF;
defparam sp_inst_14.INIT_RAM_39 = 256'hFFC0000000000FFFFE0000003FC3FFFFE01FFC018CFE000003FFF80000000007;
defparam sp_inst_14.INIT_RAM_3A = 256'hE0001FFF000003FF8C000000003FDFFE01E0003F003FFFE003F8001FFF000003;
defparam sp_inst_14.INIT_RAM_3B = 256'h00FC001FFFF00000311F3F000001FFFE000000007F0FFE03F0007E003FFFE000;
defparam sp_inst_14.INIT_RAM_3C = 256'h0000FFC3F01FF800F0001FFFF00000039DFF8000001FFF7C000000FF0FFC0FF0;
defparam sp_inst_14.INIT_RAM_3D = 256'h0000000FFFFFC0067EFFE0003FF000E0001FFFFC000007BF3F8000000FFFFF00;
defparam sp_inst_14.INIT_RAM_3E = 256'h83FF8006737FC400000007FFFC1006C4FFF0003FE001E0000FFFFF000603FF80;
defparam sp_inst_14.INIT_RAM_3F = 256'h79FF8001C03FE001FF0000F67FDE00000003FFFE031800FFF838FF8001C01FE3;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[29:0],sp_inst_15_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b00;
defparam sp_inst_15.BIT_WIDTH = 2;
defparam sp_inst_15.BLK_SEL = 3'b010;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h13C4647A4A885770821160F8E43FBF0C2C2E890085362A75C8A26C72A8467319;
defparam sp_inst_15.INIT_RAM_01 = 256'hB3EA94A758E609589829F44A79223C59DFBC3FE9AFFFD52CA7F854C41AF17AED;
defparam sp_inst_15.INIT_RAM_02 = 256'hAAA5B3652B5A99FA5E541AAC7FC4433A56AD0D57FC85B8C37671E2ABBF2EA33D;
defparam sp_inst_15.INIT_RAM_03 = 256'h4FD406C00CFE95864EABF014283DFABE16226451D27A04010FF9B66914878AFC;
defparam sp_inst_15.INIT_RAM_04 = 256'h37DE3CCE6F45CBBA8C5C6AC0657AB0002EE5F1950BF464AAAA61767C2C99263B;
defparam sp_inst_15.INIT_RAM_05 = 256'h672A51BED5CBEA8868C80686B5B6CC4962C3D6C1428DB03E006CB50CFA2FCCE4;
defparam sp_inst_15.INIT_RAM_06 = 256'h1F32331C614E156112591B3BE62C8E92AC4A721BA4D2F20CB696F42A69002EE2;
defparam sp_inst_15.INIT_RAM_07 = 256'hA158451C21BC5552EC396AA959ECD8802470378CFC48CA4B520A1BD9934EC913;
defparam sp_inst_15.INIT_RAM_08 = 256'hA470C24BC932C75459A8389FF7B86D2658F7BCFF1607E6504B7C759A83E8BD04;
defparam sp_inst_15.INIT_RAM_09 = 256'hEFFF40169537900CF8A96D3FA9A413BE5E3925BA4BCB10AAD8BE03A0D9E6C903;
defparam sp_inst_15.INIT_RAM_0A = 256'h678EC4781B1D21540E694F9BF7F8A96C07656156A7B8EFB4A4C706C893C54127;
defparam sp_inst_15.INIT_RAM_0B = 256'h65BAC4A2F436F04ADC9BF3F5BA0C3FFC001B078A513EAA0900B39E29DA141791;
defparam sp_inst_15.INIT_RAM_0C = 256'h48884776394D1D7D40FE98DB0445F90AF20E3DE2CA905400E9003753AF20FC4D;
defparam sp_inst_15.INIT_RAM_0D = 256'hDD2FF153E3A214E493AA56B0AACD80CCF37F66EE3530FF2F87DC710E4000555A;
defparam sp_inst_15.INIT_RAM_0E = 256'hD7FF729DEECE12D0277B414095556C3C9A920DFFAD49387A52269BE9FFED1EC3;
defparam sp_inst_15.INIT_RAM_0F = 256'h4C3A6C46B05FC37093102A193F23255DF4BF6D521A483A9BFAA5B374151842FC;
defparam sp_inst_15.INIT_RAM_10 = 256'h200675532CF100FE83CA804D86D0845547AFC9D9D295EF8F4FF1AA5A331A2AEF;
defparam sp_inst_15.INIT_RAM_11 = 256'h712C9E7518FE9FB6AAAFADA6A6C41ED4FD7F043BEDDB7C11C8D26C0CBB771F86;
defparam sp_inst_15.INIT_RAM_12 = 256'h6754625716C57B126FE6304EA19EBF13AE00BA7B0DD0C5EA9A3EECC398E055EB;
defparam sp_inst_15.INIT_RAM_13 = 256'h25BAABD1983BE216DF7A14CDCF55105EDBD87F2AD4016BF0615B6368A09A2CFE;
defparam sp_inst_15.INIT_RAM_14 = 256'hE15E6FDF6AAF8C1C7288235D7062C4D2B381915402AE6EC72D2A0490667566C0;
defparam sp_inst_15.INIT_RAM_15 = 256'hE5647A541B317C206F580F1E211045B62DEDBDF243FF34D236C1A480FBFE9F3F;
defparam sp_inst_15.INIT_RAM_16 = 256'h72A47B874E37A73A18E532A157AE548C750656CE3DC54D160F7548B34CBCA918;
defparam sp_inst_15.INIT_RAM_17 = 256'hF8CB76F32F939D04EA76A397F85205D0555513AFBFD38C8EDB8998431296E279;
defparam sp_inst_15.INIT_RAM_18 = 256'h911B8FC6BF948CDA067B1CCDBC96D52068461B00E5B3053A687FED01C1D4643D;
defparam sp_inst_15.INIT_RAM_19 = 256'h39562644653E74A23A94DAF1362F018C0F3267357D6231A697613570009541AA;
defparam sp_inst_15.INIT_RAM_1A = 256'h9463DE62598505BA6151F34651BCA10DCC3D0E846EF68CF1522849FE4C9EEB85;
defparam sp_inst_15.INIT_RAM_1B = 256'h107DF7313B3D026BD7069E3F3B3C00F4F4F4BD02E3993FAB33D7C97A0BDC67F3;
defparam sp_inst_15.INIT_RAM_1C = 256'h3974A274B5A2D313DAD7681C30F033467D613C0BAF251847F096516F569640DC;
defparam sp_inst_15.INIT_RAM_1D = 256'h30FD28DA4A3AF1E6416A063C56C440ADB2E28929E76AFACE9E8B0AD7F125421B;
defparam sp_inst_15.INIT_RAM_1E = 256'h1309FA1AE1FE220FEF54030882107B3270760BDA522790AC32721729E90C96C3;
defparam sp_inst_15.INIT_RAM_1F = 256'h7936373D644AC1DC6216EBA9C99F6CB3246D1C7CABE50169050DEF3E69344FC0;
defparam sp_inst_15.INIT_RAM_20 = 256'h025CD1AA955504049BFAD736740B03AA8D6F593757AD8735C29AD91371EF900D;
defparam sp_inst_15.INIT_RAM_21 = 256'h5FF5A761BBEECD89B19980B889A78B5A9FADD976FFC12A3E425DE9C5BD20A748;
defparam sp_inst_15.INIT_RAM_22 = 256'h8A6B372D431405138319D4A0A04E30B575C639550402DA3EB13B1AA54D4E156A;
defparam sp_inst_15.INIT_RAM_23 = 256'h9B6AA55681B34960B618B597E4059B2CAAEAD0BFEDDB3FDA47D970B23BCC140B;
defparam sp_inst_15.INIT_RAM_24 = 256'hAAD494793FB813E6E643B9BC95E8E04069D3F4E1F86E1C3027E531C871A03F71;
defparam sp_inst_15.INIT_RAM_25 = 256'hE98BF22A477497A07C595E3DDF8F44FCE4068723998BFFDF537EA0906B2AF295;
defparam sp_inst_15.INIT_RAM_26 = 256'h614D4CCA9CD34BC33ED24E4C5A6F6E07383631F19FD1E0749C549EFA752CCA56;
defparam sp_inst_15.INIT_RAM_27 = 256'h800A65172D4BD1AA80525AA79BB99E0726FE6F181F007B954C8DBDEA22952005;
defparam sp_inst_15.INIT_RAM_28 = 256'h486D2E4077F9A4AEF025758EC405D496950C1CD5B4ABED202C8DD4040B22D824;
defparam sp_inst_15.INIT_RAM_29 = 256'h80AA5FB69655688041B2EA3FE5E0AB03849EA90A2CFA5478AF6042B81A822B37;
defparam sp_inst_15.INIT_RAM_2A = 256'hC26B9C85AA553758B4DABE72A34A2CAE3A06AEC2BD4D2581E1F81901757C7234;
defparam sp_inst_15.INIT_RAM_2B = 256'h82678AD7E864683FD900A6662BA466D4127C0A21AE147E85ADBF583A1285C618;
defparam sp_inst_15.INIT_RAM_2C = 256'hFDF1AADD011A30D57B596E0D7B9529A7EE2BE064CCF42A9EA19DF4528EB5E915;
defparam sp_inst_15.INIT_RAM_2D = 256'hFC55F9302BCAE2956666DD7B3768C84A4EB01AA5C9998900002E15704E9CA968;
defparam sp_inst_15.INIT_RAM_2E = 256'h6A5654A24E4100EC78299A9F11C4BDD8EC7640034B400C1579618B0D3CDABE33;
defparam sp_inst_15.INIT_RAM_2F = 256'hE8933A76ED423FEB37CA5F2E364DC3322163C81C64F613A82BB521E32C83A6F2;
defparam sp_inst_15.INIT_RAM_30 = 256'hAD8D8BABEBF84AB962FDCE2A6FD2AAAAC73DF91D0D17DDA3BF4E6AA7A8C9CF1A;
defparam sp_inst_15.INIT_RAM_31 = 256'hFD0D6C73675675B5780DAC70C312C68651E076B7A7DC2CFD93318D11F331CB93;
defparam sp_inst_15.INIT_RAM_32 = 256'hDD1F70D19E2705E8A921A450F7925D15C2A4761874273C596C29ADF305004C02;
defparam sp_inst_15.INIT_RAM_33 = 256'h47AAEAA6E20208DE5CD2600F2FB4CE0D810B0573C36C48B3022914F3074E8A9D;
defparam sp_inst_15.INIT_RAM_34 = 256'h6D533CE9387FDD51C4FE97F3C563D3AD514678C4AFB5CD6B2325EF0AD4986EF0;
defparam sp_inst_15.INIT_RAM_35 = 256'h2E64CBF06D6F600DC3074F53A990BAE030F1C9622C9201681D43858FC20E3507;
defparam sp_inst_15.INIT_RAM_36 = 256'hED29BC374B302150A22A870D0B1C4F00C6158A0F363BF014B38FEC94D701DCDC;
defparam sp_inst_15.INIT_RAM_37 = 256'h79EBB0000FC053F011774E23F9DBCF618141EE95DAF622CE984838F41D66FFAC;
defparam sp_inst_15.INIT_RAM_38 = 256'h0A41E10D229D785D15A3EBECAA80D35A78AC733E5FE91395844921CB2B4275D8;
defparam sp_inst_15.INIT_RAM_39 = 256'hA386FFEA5A5584987F5025D34AA1A203ABC14FFFC513351F8314F2962B485CCB;
defparam sp_inst_15.INIT_RAM_3A = 256'hF140BE813BD7D7268C38253406CAD5BAA7A4A3F276A0E867CD4491538AC77CEA;
defparam sp_inst_15.INIT_RAM_3B = 256'h8A385ED3423A4AFE01AF395B50167EBF0000001685E8F383D683BE76F0C66F58;
defparam sp_inst_15.INIT_RAM_3C = 256'h1405B5C716A2896D6C57C77B98E768C3000F0D6F9C6E304929BA81AE15694947;
defparam sp_inst_15.INIT_RAM_3D = 256'h0EA90D49385E23B741F3985D9DB8FD72198EC8593ACF55BFE96A43FF5E6F0015;
defparam sp_inst_15.INIT_RAM_3E = 256'hA54A3FFFAAF0AABF50FE5EB040151541B5C2FB472149FF51F8000898561653AC;
defparam sp_inst_15.INIT_RAM_3F = 256'h132296A6B9A2BCB97C22FDD2FE58FEA7E5333A2B2825CF82AACE7B1B7FD6CB0E;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[29:0],sp_inst_16_dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b00;
defparam sp_inst_16.BIT_WIDTH = 2;
defparam sp_inst_16.BLK_SEL = 3'b010;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'hCD6A0005D5FDFF050054EA555540006BEBEBC000FFF33FF0C13E428076BEE83A;
defparam sp_inst_16.INIT_RAM_01 = 256'hF3FFFFB30103FFF90140A2ABFFE99500154FEAAAAAAC0EABDFFF9E6AAAAFF150;
defparam sp_inst_16.INIT_RAM_02 = 256'hAAAAAEAC4EAAEFFF9EAAAAABF150FE5075C89126ABC0F1143E45540000555AEB;
defparam sp_inst_16.INIT_RAM_03 = 256'h200BFFC00100035550000555AAACFFFF03F3F154A9540154B2FFEAFFFE03153A;
defparam sp_inst_16.INIT_RAM_04 = 256'hEFC03F50007DEFDE5163AF4154EAAFFFFFAC03AAEFFF93AAAAAF05417BB5A94D;
defparam sp_inst_16.INIT_RAM_05 = 256'h03EA8AAA53BFAABC5516A3141AA70D5EF014001403A505405556FEBCFF0010FF;
defparam sp_inst_16.INIT_RAM_06 = 256'h4F0433E50550555AFEAAFF05533BFAB014A4047CFD96F39732D154EAFFFFFFAF;
defparam sp_inst_16.INIT_RAM_07 = 256'h46A4F187EA9EE7A550EAFFFFFFABC0FFAC053EBCABC164156453C56A3050C1A9;
defparam sp_inst_16.INIT_RAM_08 = 256'hAAAFBF1564045557AB1BFBC005AA4FF0009401005555AAAABF069EFBFEB12B82;
defparam sp_inst_16.INIT_RAM_09 = 256'h00005555AA9AAFB15ECFEBF012825A90C7E6A969B4E593AABC005400C0FFABFE;
defparam sp_inst_16.INIT_RAM_0A = 256'hA964A5403AFC5AAAA5555000FEAAAAAB0055540019553AA2F7BF556503C01794;
defparam sp_inst_16.INIT_RAM_0B = 256'h0000501A952A03FAC153AF03FEA540015555BEB9AF9D4A653FAE0F0E7EA462AA;
defparam sp_inst_16.INIT_RAM_0C = 256'h6D3BB0DB3C5190EAB13AFC080BBF96F7944FEBC56AAAAAAA555543FEAAF00150;
defparam sp_inst_16.INIT_RAM_0D = 256'hBC555AA9A95AAA55540000050010C01179ACAF89AFECFF000EBC3EA555555555;
defparam sp_inst_16.INIT_RAM_0E = 256'h8BE3AEB253BC54FF3E9555555555AB00C000013C553A053FEDB4DE6A969E903E;
defparam sp_inst_16.INIT_RAM_0F = 256'h0C3FC64F05538A658AFFEA7A406E0550F1559005AAA540000000F30500569396;
defparam sp_inst_16.INIT_RAM_10 = 256'h40005AA94FAF00FFC3C015516A4E6DA4F98564ABC553AAA55005555563F15550;
defparam sp_inst_16.INIT_RAM_11 = 256'h04EBC0053A55500555559700064C0FFAB14101402F256DAA50A9016C543EAB15;
defparam sp_inst_16.INIT_RAM_12 = 256'h94ED59D66ABFE954001194FAAFFC005401AA4EAF50FFC0FF157AB2B8E6C3AA84;
defparam sp_inst_16.INIT_RAM_13 = 256'h93C554FFFC3F1A896B6F8ABA6AB003ABD9014E955555555AA98530ED14E6FC01;
defparam sp_inst_16.INIT_RAM_14 = 256'hC4E5555055556BF244AC5294F19315EAB4F7155AA90000114FEAFFAC54053C6A;
defparam sp_inst_16.INIT_RAM_15 = 256'h014540000041EBEAAAADA2B17CAAA4195501EBF06FE3EA8BD3AAEA6FA96C2FD3;
defparam sp_inst_16.INIT_RAM_16 = 256'h6AAC5AAA8A9D0E9B4E6A9AB3D9B9FD4A6FFD5565ACFCD525E9546057B9B6A75B;
defparam sp_inst_16.INIT_RAM_17 = 256'h5515A12C003966AEBC79612D4AC555000000000B96A9A6BC498656AAA450546F;
defparam sp_inst_16.INIT_RAM_18 = 256'h000BA56AAAAD516AAA95A0114C7E7BEC5506F8EAF965A795AABD6B1B9E9BBE5F;
defparam sp_inst_16.INIT_RAM_19 = 256'h6E39FE8A1896AC7CEAADB35339BD1A51BF0417EA269B54E97EC4C43C55000000;
defparam sp_inst_16.INIT_RAM_1A = 256'h853EB9AB64A9A74F57FB040000010007BA96FAA856A9165AA70150150FB15550;
defparam sp_inst_16.INIT_RAM_1B = 256'hAA97F043AF06A7FFC3FFFA1440411A3FB0B4B3AAC41BDEAA0540CEB390651C3E;
defparam sp_inst_16.INIT_RAM_1C = 256'h3EAAFEAC6E2A443014C3E556D6C39B505A4EEB95AD7793FB050000000006BFA6;
defparam sp_inst_16.INIT_RAM_1D = 256'h9506B59C6C41050000000042AABC69D15AA9BFF152AAAABAA8503B1405400004;
defparam sp_inst_16.INIT_RAM_1E = 256'h03FC4EAAAAAAB542D9B15450E6F0945A4EA98B8A947A3FF4AE45BD61FA252DF1;
defparam sp_inst_16.INIT_RAM_1F = 256'h97A72C302ABAA5655C25D46734886559AC1092C5000000000052E5B6FF8EA56A;
defparam sp_inst_16.INIT_RAM_20 = 256'h556E000000000052394FFE91EAAAFEAC4AAAAA9A146BF8DB140E92EF9ABCF8E6;
defparam sp_inst_16.INIT_RAM_21 = 256'hAAAC55FFEA9EBC0F9698EB0FFD89B9D4A6F2EAAA556A960EB19F1535A6EC1E0C;
defparam sp_inst_16.INIT_RAM_22 = 256'h155443E57D6256250314E7C69500D545401540000051FE9FEE56AAAAA6B27AAA;
defparam sp_inst_16.INIT_RAM_23 = 256'h52400000CE98151B6EABAFD8AAAAAAF21BFFBF8A6580256CBFE655D9D622AAB1;
defparam sp_inst_16.INIT_RAM_24 = 256'hE3FA83FF39BEAC49561EEABBAB155556550396AADADCAEF18F0EF515E456AC5A;
defparam sp_inst_16.INIT_RAM_25 = 256'hE6FA6C438A7FA13D5867ABEABFFAF9E500008EB3FC11696AEBA2A1EAAA141FFF;
defparam sp_inst_16.INIT_RAM_26 = 256'h7FFAA7F96BAA868AC503A851BFFF4FEBBE2AF3AFAEDFA65715EAC0F1559F1555;
defparam sp_inst_16.INIT_RAM_27 = 256'h6C3ABEBE09A0D2AB53AF55396C555EAAFAC5EDA4B51605B940C0FFAA940E4000;
defparam sp_inst_16.INIT_RAM_28 = 256'h654254C24401404BFE403FCF50004FFEA6E66A6C7CAA9590C650BFF90EA7FA7A;
defparam sp_inst_16.INIT_RAM_29 = 256'h33DACAA1003C550EC6FBF9DFFE3FAAFEAB9075D976AD3AAAA1DAAAC6A7AA1459;
defparam sp_inst_16.INIT_RAM_2A = 256'h1305AA47AAAA99754E6C552C3F01C626452540175C1E956A54FF9000443FE5EA;
defparam sp_inst_16.INIT_RAM_2B = 256'h0404A26A56AAAA7950003454FAFF1AA5AE8A80A58A9658B794BEF89A9556BEAA;
defparam sp_inst_16.INIT_RAM_2C = 256'h05C9526AAAF993FFC9BE998546AAD4D15611AAAA66D7C4965A29E22D2717328E;
defparam sp_inst_16.INIT_RAM_2D = 256'h56AA576010AD5A7DF4A1BAA2701990673F5BAAAA6A49500063156A9AFA76AAB1;
defparam sp_inst_16.INIT_RAM_2E = 256'hAAAAAA4D500014FBFC3F990EAAA810525679AAA94FFE62957B8E508D6C35667B;
defparam sp_inst_16.INIT_RAM_2F = 256'h56A98AAD96597E2995F6559156255A999A0404C66A7B9313AFEAA8C47A056DD5;
defparam sp_inst_16.INIT_RAM_30 = 256'h0E869679B0EBFAAC5D9E85DBF5DBAAAA697A0001394FF5AA7797AAA9B11665A4;
defparam sp_inst_16.INIT_RAM_31 = 256'h0001279A8DC1ECA39BAA015A69A9496AFF2DB99AF7AA985EB5896984181E1284;
defparam sp_inst_16.INIT_RAM_32 = 256'hE54FDEA53DF5FFFAAE73EBF1066BFAAC1A7AAFEBEAAFEB15297C5524AAAAA539;
defparam sp_inst_16.INIT_RAM_33 = 256'hF9BEAAAAAF9EA4B15C345AA59395100127FFF98935EAA6AF55AAAA596897A6C3;
defparam sp_inst_16.INIT_RAM_34 = 256'hF6505996AAAD16AA6A55554D6BEE553E7F90F6FFF3F514EAAF555F4AABFAB12B;
defparam sp_inst_16.INIT_RAM_35 = 256'h9FCE8FF0F83BC5BA7E7FFAFE9DEFAABEEFAFBAC2F27A13D901540E5014015153;
defparam sp_inst_16.INIT_RAM_36 = 256'hABEBFA1755A9AFFFA9401401595CF2E452B13AD75A955AAA5950A8EA6BFB801A;
defparam sp_inst_16.INIT_RAM_37 = 256'hE70D5AAAA56AA95ADE4A96A0ED7E49AEB3FA0C510F2EDC79BFABF0AFABEAAAAB;
defparam sp_inst_16.INIT_RAM_38 = 256'h4F0EBDAE967FEBFAD2AAAAABAAAA73F9FFAE854255555400150144CCC0A59F96;
defparam sp_inst_16.INIT_RAM_39 = 256'hFEB600000000150142FC3FD8B9D25918556AA5556AA9952469AA04FA213B9FDB;
defparam sp_inst_16.INIT_RAM_3A = 256'h5AAA556A95525595551C8F47E581EF02AE0D18FAEAAC7BEABABFAAA9FABFABFA;
defparam sp_inst_16.INIT_RAM_3B = 256'hD8FBA6B5FE9BFAAAAAAAEAAAFFFFAAAA0000000015010654C067DBA164665556;
defparam sp_inst_16.INIT_RAM_3C = 256'h00000500428469012BEB455569A1AA69AAA5A55521557773C1F4EA5BFAF1E19A;
defparam sp_inst_16.INIT_RAM_3D = 256'hA555535509A7AA5D0EDA4BE8176F4AEAFC12BABFEABAAAAAAAAAFEAAFAAA0000;
defparam sp_inst_16.INIT_RAM_3E = 256'hAACEEAAAAAAFAAAAFFAAFAAF00000000050005A09E6F3EF115A69CB41A95A956;
defparam sp_inst_16.INIT_RAM_3F = 256'h55A1468C7F039A5A47FDE86955565554506807990F3A3E9E9783804C2BFF153F;

SP sp_inst_17 (
    .DO({sp_inst_17_dout_w[29:0],sp_inst_17_dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]})
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b00;
defparam sp_inst_17.BIT_WIDTH = 2;
defparam sp_inst_17.BLK_SEL = 3'b010;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'hB8AAA8A89D28805FFD5F2A20A22A0A00A20897DF8AAC402D9F400280ADFD77EA;
defparam sp_inst_17.INIT_RAM_01 = 256'h8C0808267FDC2A808A882DD77F7F7F7DF5F882200203F02A37FFF8002A8285D7;
defparam sp_inst_17.INIT_RAM_02 = 256'h28000A03FA8A15FD50220022A777888F48B89FCA80370D5D42A88A82AA8AA2A0;
defparam sp_inst_17.INIT_RAM_03 = 256'hFDDA2097F55D548A0828A228AA0B082AD62E8575AA880008AFFFF7FDF55477C2;
defparam sp_inst_17.INIT_RAM_04 = 256'h28BDCAA0A088BD5A882FDFDF558A2820A02B7C8A37FFFC208280DDD5C2057D52;
defparam sp_inst_17.INIT_RAM_05 = 256'h56A037FD7CA0A8A3FF777CFD75FC5378AD7F77775682082A2080A8098AF75F20;
defparam sp_inst_17.INIT_RAM_06 = 256'hD2FFCE888A800A8A80A222DD7C60AA85DD0A2280F588A4A2CD77DF2828822008;
defparam sp_inst_17.INIT_RAM_07 = 256'hAA80741F5F702A55D722822A28023F8A835FE28B8A355D775D7E35FF65DDB5F5;
defparam sp_inst_17.INIT_RAM_08 = 256'h2208A8D777FF5FFEAA55DCB7D5FF788FD7A808AA8A2228222AFDD208A00D7CBC;
defparam sp_inst_17.INIT_RAM_09 = 256'h88280808A2000825FA9008AF7C948A2AD0DF5755A0B57EA0095FD57517808028;
defparam sp_inst_17.INIT_RAM_0A = 256'hD7F5803762A9FF5557D55FD728A8088AF5755FFDDD7D4A2774887DF776155C88;
defparam sp_inst_17.INIT_RAM_0B = 256'hDD5F5557D7EA5E8A15DC8A74A0A2800AA2000A28080BD8DDC288FAF0288A675D;
defparam sp_inst_17.INIT_RAM_0C = 256'h8368A700CB755F800F6021FA7DFDF5F60A98A81F7FF75FF77FDF5E22880D5DFD;
defparam sp_inst_17.INIT_RAM_0D = 256'h895F555F77575757DF575DDF57FF3757EA83D558828388DF5AA340A8A200A082;
defparam sp_inst_17.INIT_RAM_0E = 256'hBD5C00077C83DD02CAA8282A00882A5DBF7D7DC35F6AF5E2AB4A1777D5788880;
defparam sp_inst_17.INIT_RAM_0F = 256'h7B68BFF2FF741D62B557DD60A020F5DD87D775D7F555DFD757F7AC5FFF75DE22;
defparam sp_inst_17.INIT_RAM_10 = 256'h75DDFF5FD002F500341F7777F572895F881D77A01D5E0AA0A00228080EADDF5D;
defparam sp_inst_17.INIT_RAM_11 = 256'hDD2017776A082828A28880D5FD79FA288FD75F5FF76029D7FD0A28837D4088F5;
defparam sp_inst_17.INIT_RAM_12 = 256'hDD8B578A2200220228AFFF008281FD7DFF5DF228D528952055C88D7F08BEAA15;
defparam sp_inst_17.INIT_RAM_13 = 256'h7E37D7882BCA7F7088D550AA002FF4A09D7550A8828A22022815450355AA09D7;
defparam sp_inst_17.INIT_RAM_14 = 256'h958AA208A22802AFF7A3F48B257EFD8A2F27800AA0A0A287588A200B7F554957;
defparam sp_inst_17.INIT_RAM_15 = 256'h22AA288A80AD88A20829548763F55577DFFF202577F400B7F6A828AA20A3DF7C;
defparam sp_inst_17.INIT_RAM_16 = 256'hCA8B7DFFDA2BD080F888202EBFF70BF028022A000381356800A17DD6AB60A25D;
defparam sp_inst_17.INIT_RAM_17 = 256'h2AA8A561DF4882A0A168A741F83D0AA0A8A2AA82288808A35897DFDF7F5FDDF7;
defparam sp_inst_17.INIT_RAM_18 = 256'hA8AA08A80089D55F7DD7FDDD5B7DEAA9755DFF8828ADD60A88202A5552962A28;
defparam sp_inst_17.INIT_RAM_19 = 256'h7FC0009D5580A1770029D456E2AA2202A8FD7608C0AA570A8A1F3FE1822A8A8A;
defparam sp_inst_17.INIT_RAM_1A = 256'hB74AA2807FA20050DC080088A2A80A0A8002A82BFDDD77F5D47F7575D2AFD755;
defparam sp_inst_17.INIT_RAM_1B = 256'h808207DCAADD7EA21EAA00FDF75D5DE00DA72488BFFFD0A05FFF322402A2814A;
defparam sp_inst_17.INIT_RAM_1C = 256'h6AA880237548354F7D96A0AA803CAA5D5A088A88A36F76A208802A808A282A0A;
defparam sp_inst_17.INIT_RAM_1D = 256'hA02A0DBF2BF7000A82202AA8A20B7F22200A008D7600A22A0355E85FF7FDFF75;
defparam sp_inst_17.INIT_RAM_1E = 256'h74A9502228AA255FF0077757008F2282F0A8B5F8B5CA4082822A28AD2A77EB0C;
defparam sp_inst_17.INIT_RAM_1F = 256'h827463C5E20822A289EA1D5C473200AA09D48ABF2202022A8200AAAD7FD8A8A8;
defparam sp_inst_17.INIT_RAM_20 = 256'h8A2082008A0A08A8683D5DF6A0A0A2A9D002222055FFDF02F7F282208A235720;
defparam sp_inst_17.INIT_RAM_21 = 256'h8223F7FFD770A9FA0A29027829F08ABD082728AAA8A80AF08578FDCA08A3FA5B;
defparam sp_inst_17.INIT_RAM_22 = 256'hD77FD4280205DD6DD6753C37D775800BAA8A0A800028809D7D562282A82FC808;
defparam sp_inst_17.INIT_RAM_23 = 256'hD688220AB81D5F5E82080A9D800202875D55DF58809FE2A30A8288BD0AD402AD;
defparam sp_inst_17.INIT_RAM_24 = 256'h5400BE82EA880378AA8363E028FDF7F7775620801D8B588FD25AA57DA008AB77;
defparam sp_inst_17.INIT_RAM_25 = 256'h880201F4BD68A7E0835CAAA87FFFD5A2AA02300CABF6AA20AA7E072A205F7D7F;
defparam sp_inst_17.INIT_RAM_26 = 256'h82A8202882221FF83DFC0355D7DFF88A7D688EA8ABF2A808D588978DDFF87D7F;
defparam sp_inst_17.INIT_RAM_27 = 256'hA968A0A850881488DC005F40A3D7D022803529FF8FD680229737D57777720820;
defparam sp_inst_17.INIT_RAM_28 = 256'hD775DD368A22155AF5DDCA32888A92A0A88028A37F0ABD771D7D7DD7D0055DE8;
defparam sp_inst_17.INIT_RAM_29 = 256'hAE97520FDF49FDF03DF4A0BF57600A8A808885A3688968AA8F2A089F7E8A7D57;
defparam sp_inst_17.INIT_RAM_2A = 256'h2DD528BC2A28A2A55089D563C8DF95CA7568A220A9D87DFF55A80A821FE88A82;
defparam sp_inst_17.INIT_RAM_2B = 256'h8889841CD7F5FD4800A8A7F702A8FFDFA09D7D0D728A89DEAB7DDFAA82802AA2;
defparam sp_inst_17.INIT_RAM_2C = 256'h7D1DD48202A885DD7A2AA152AA82239E2074800820961D20D7C32D4960FE45D0;
defparam sp_inst_17.INIT_RAM_2D = 256'h0082806A2FABF7C32F0F022D4777A282EAD27D777DFA82008477F75557E022AF;
defparam sp_inst_17.INIT_RAM_2E = 256'hF7D5F5D2A82A872801E0B7D8820BD7D5DDE2A822B77D40A2877088122360A84A;
defparam sp_inst_17.INIT_RAM_2F = 256'hA0AA155D0A2A7D62AA80202A2AC08220A0D8B797F7C25C762AA8F53F40086B8F;
defparam sp_inst_17.INIT_RAM_30 = 256'hFA1D5FCA85022A838BDA3FA8AD3E55F77FEA80280F72A0A8043C28A82577757F;
defparam sp_inst_17.INIT_RAM_31 = 256'h88A8A628103F01768800555F5DD5FAA2087500A3D4208388088AA977DFDDD495;
defparam sp_inst_17.INIT_RAM_32 = 256'h2AB7FA0220A00AA82B6C2A2DD5C022815F6282088A2AAA75C963F7FD75F5D7C0;
defparam sp_inst_17.INIT_RAM_33 = 256'h082200280A895FADDB49555F54AA2288A68222374F288288F5FDFFDFF5882A16;
defparam sp_inst_17.INIT_RAM_34 = 256'hA0577D80A20377F7D55D7D5082A0087FC88A22A22C822920A257F2D8228AA7E8;
defparam sp_inst_17.INIT_RAM_35 = 256'hA2B2300FA142BD7D5E202A88090A0A0200288A34856AFCA1DDD572A228828DDC;
defparam sp_inst_17.INIT_RAM_36 = 256'h0888AAD40AAD28228880A202A17B257FFC0FE0167D75DD7D7FFD890800FD7D20;
defparam sp_inst_17.INIT_RAM_37 = 256'h1471775F7F75DDFFD0A80AAF7222B888A62AF155D0D5D70200A82D28880AA882;
defparam sp_inst_17.INIT_RAM_38 = 256'hD0F2AA15D42A88883C028A2080A00CA22009FDD60280022AAA20031B1DD52A3C;
defparam sp_inst_17.INIT_RAM_39 = 256'h208A8A200AA0AAA28A0342158034FFD5F77DD7FF77D5FDC08002FAAACDE0A2B2;
defparam sp_inst_17.INIT_RAM_3A = 256'h57DFF7FDF77EA000214B3D5C0015885E0A2B58AA80A3E2828088A880AAAAA800;
defparam sp_inst_17.INIT_RAM_3B = 256'h9A08228FA08AA082A2280228A8008A0AAA02A028A82008D7BDDC08A7777DF7FD;
defparam sp_inst_17.INIT_RAM_3C = 256'h20220A2A8A7DD5FD4008FDDDF5A577D5F7D5D77FC008AC861D5500A2A22D8F80;
defparam sp_inst_17.INIT_RAM_3D = 256'h5F7576A07282A850B7A2D8ABD40A500801F4A82822882A2AA28AAA2882222828;
defparam sp_inst_17.INIT_RAM_3E = 256'h28902A2A808202A080AA0AA208202028A28A02D75AD8680DD75DDBFF5FDFDF7D;
defparam sp_inst_17.INIT_RAM_3F = 256'h2ADDFF5B4A7CB55F57FF295757555F5D75C940A272C0F7D03496F7D1622ADD42;

SP sp_inst_18 (
    .DO({sp_inst_18_dout_w[29:0],sp_inst_18_dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]})
);

defparam sp_inst_18.READ_MODE = 1'b0;
defparam sp_inst_18.WRITE_MODE = 2'b00;
defparam sp_inst_18.BIT_WIDTH = 2;
defparam sp_inst_18.BLK_SEL = 3'b010;
defparam sp_inst_18.RESET_MODE = "SYNC";
defparam sp_inst_18.INIT_RAM_00 = 256'hF7B4F952354CB2152867A3EB92956A0C37D4E3A5EA48251FB6F16C4786AC8B24;
defparam sp_inst_18.INIT_RAM_01 = 256'h2A503E3C4648F3A8583AD2E3BFDDE75A8B87FF3FEB5B9D6F2FF8F87EAFFF1D9D;
defparam sp_inst_18.INIT_RAM_02 = 256'h5BFFEB06E26ACD65BDBDB0EF12B44D4BFBC9F8235B6F1D1A8A7198C56F2ABEEB;
defparam sp_inst_18.INIT_RAM_03 = 256'hA6E0F16A1105E58634F1B0552F36A5546CB7643B88CB495298FEBBBF6F44252C;
defparam sp_inst_18.INIT_RAM_04 = 256'h47C5E6136056FFBA38AC2B7FC2FFAC050546F8A57EA387FEC3B1863C2F3D6651;
defparam sp_inst_18.INIT_RAM_05 = 256'h6DEA2F10D8C50FB617BDAD11A5BB1601C700DB18428D5540F1767D355073D24E;
defparam sp_inst_18.INIT_RAM_06 = 256'hD074FED81555BC77D90DB046578B24D1169EB62CF78D220C23F161EC00C3F00C;
defparam sp_inst_18.INIT_RAM_07 = 256'hA56C80CBE1BFF1F8A13EC30396F8DE0FA185E7D50F1C6141577E1BD955B008BE;
defparam sp_inst_18.INIT_RAM_08 = 256'h3EF901851009733759BDA9FCFDC8137B0263A5062C5CED77DC7796057E781204;
defparam sp_inst_18.INIT_RAM_09 = 256'hA696ABC63FF49FE5B8AE188F3964DDEF99B97AE4A711166F6DD43B5CE355A8F3;
defparam sp_inst_18.INIT_RAM_0A = 256'hBB83B3E3CF07B1BF69673BEA93C30FAA07551DBC58C243A51142E8BB27F1F9E4;
defparam sp_inst_18.INIT_RAM_0B = 256'h25CFA8ABC7E7DE05185603F6660CFAABAF1B58264C93BAC56A19472384140791;
defparam sp_inst_18.INIT_RAM_0C = 256'h48DEDB8887D4C994D39932D83435F909A945E886EAA96AA9400F483E6B160C09;
defparam sp_inst_18.INIT_RAM_0D = 256'h877F3AA39406A9530FFFABC0FECDC0CF5730D16DCC33507ED7D1710E3FFCF01A;
defparam sp_inst_18.INIT_RAM_0E = 256'h82F63386806612EA377B3C3C55161838D4339BF0B0509D64A7779BD8FF84C55E;
defparam sp_inst_18.INIT_RAM_0F = 256'hB42B1DFBC04510B442CED5F3EBAA75139614B4C86E54ABFFAAA9C04465F2E6FD;
defparam sp_inst_18.INIT_RAM_10 = 256'h256BD95634EAF000C41AC3D61F2599B1988F1386DD963F8F3FF1AAAB3300CF36;
defparam sp_inst_18.INIT_RAM_11 = 256'h981687D1580F8AA2AFC1B29F3AC9AD851299F31FDCDB6BCF62B75882A75254B1;
defparam sp_inst_18.INIT_RAM_12 = 256'h4E37AD51F0A3D1FC5B56ECFFFFF2C6F95B0786B1BE2BDA7F844F0154F0A6A9DC;
defparam sp_inst_18.INIT_RAM_13 = 256'h489D16EBED4C766CDC8F2679CF94C14B8CD27F3F93FCAF1AC893C8AC9F5F7B52;
defparam sp_inst_18.INIT_RAM_14 = 256'hA2635A8A6F067B90DCDB7E6268F28F71EA8F0C0E585E5A3620FF434ABBDFCE06;
defparam sp_inst_18.INIT_RAM_15 = 256'h43CE81141B5C943955070F1DDE56123F84A2C34783F1E5D6B4D701EA4D264FE8;
defparam sp_inst_18.INIT_RAM_16 = 256'hCC311C73CA77B0DD6FF48BBF53A338EDBFAF3C8B81DF66774E25874AD372F952;
defparam sp_inst_18.INIT_RAM_17 = 256'h38CEB6F48E555CF42A783298BF770080015453D105ABB788D634DC576EE6ADCE;
defparam sp_inst_18.INIT_RAM_18 = 256'hE2788AB7AAA78A457B9068C86A7C9119FD42C866FECC0B1967F42C0665F0A3E4;
defparam sp_inst_18.INIT_RAM_19 = 256'h3EC63D3B6B028C714A95EA1C3A1A5AC10AF34A903D617066E26142830381006A;
defparam sp_inst_18.INIT_RAM_1A = 256'h255A9E62887305BADD4B0342006C317D1CEBF588FDB45AAA7F6B39EDAB2D3FC4;
defparam sp_inst_18.INIT_RAM_1B = 256'hB5F2FC5E6F316FC028AC99293C4C16BAA54719129DD703AC3033BABA211C66B3;
defparam sp_inst_18.INIT_RAM_1C = 256'h3E735BA7F5B385D33BD6226CF0E12B2BBDB10C065F256D410096406FA6F283C6;
defparam sp_inst_18.INIT_RAM_1D = 256'hCA4CD92F89920525005A5608F1FD8FB906F9BE860ABEAA032FB00C77F7E82E6F;
defparam sp_inst_18.INIT_RAM_1E = 256'h400172B327136FE0E0A80082B26480EBC4770BDB6937C56FF7C7572AD27A2AC0;
defparam sp_inst_18.INIT_RAM_1F = 256'h7948387BED911F66736BEB50FD807457EAD81F2BEFE400555414F5D3BFAB901B;
defparam sp_inst_18.INIT_RAM_20 = 256'h12A7E5AA505590CF367FE957391C7CB25AC3AE77A74697356ECC7D67A06EE003;
defparam sp_inst_18.INIT_RAM_21 = 256'h6F930DFBB69E65AAAAE95993856A476C4A1535C3AA5B8F4458E2DD8B99191947;
defparam sp_inst_18.INIT_RAM_22 = 256'h23A70DD04693192B3D416CE89AA62604B58134159405995F7797B6A4138E32F9;
defparam sp_inst_18.INIT_RAM_23 = 256'h561195ADA1D52E874D687923A5BFAABA93E523AFA236A06980D480AE38321780;
defparam sp_inst_18.INIT_RAM_24 = 256'hAAD49AFEACC71C12F643B337302234996E406485153A146F82ED281CFD403FB5;
defparam sp_inst_18.INIT_RAM_25 = 256'hF18578D7F5503259668D7A121F8F33AB906CFCF02AA31B2FAF2C9940F9645795;
defparam sp_inst_18.INIT_RAM_26 = 256'h5B79B84ABC66293808551A27AE7FDA027F0E5DFF70D6E184687C533536886F9B;
defparam sp_inst_18.INIT_RAM_27 = 256'hDBF0FE582D48471131F7B0AD29F7F0066597596285F8A2FDC1F6BE2ADD70205C;
defparam sp_inst_18.INIT_RAM_28 = 256'h86F3D4E9BE1D1982F0253368856B6473BB3AB9F9FCC66695CF1E1419BB72D995;
defparam sp_inst_18.INIT_RAM_29 = 256'h2AD282AA4DA68313D1B2470FE0E5BC64EDF0A90E7B505A12BFB622AF1E0C66EF;
defparam sp_inst_18.INIT_RAM_2A = 256'h4D33481A054121ADFA4E6F4BDA02E27520AC2E6AD91D25B09C93196A5673A7C8;
defparam sp_inst_18.INIT_RAM_2B = 256'h63DB1112AB1417E6DE56761735B9BD97CD1AA7C169F68E445DFC02A5D7EE6C71;
defparam sp_inst_18.INIT_RAM_2C = 256'h6A4C1681411B40EB660523AB253E0C85ED6DE5A313441497EC1D6AC329BAD340;
defparam sp_inst_18.INIT_RAM_2D = 256'h555308BA28A7BDD4D42B2E462CDBEDFDAFAA0694B0334E96DE5C8A05006D783A;
defparam sp_inst_18.INIT_RAM_2E = 256'h190603583F968474F2074462111C68960161FC05EF5B002F4F118AA1B4076845;
defparam sp_inst_18.INIT_RAM_2F = 256'h814E3487E2927C2FCF8A4AE015F32987263E67934E32B95D261FCBBC6B7955FD;
defparam sp_inst_18.INIT_RAM_30 = 256'h181606E3AB02DE8DFF19F4906C1D55050291C398F82D8710FA775569EBA9FF05;
defparam sp_inst_18.INIT_RAM_31 = 256'hC3581C855CADA6FF880EAB2CCFD2C02656B57BFBA811FBA9D3181B7DAED6D10E;
defparam sp_inst_18.INIT_RAM_32 = 256'hCD1F2C2AA593AA1591790D9F13C44CB9322090BED9B8BEA356D4F74405000AA8;
defparam sp_inst_18.INIT_RAM_33 = 256'h334E9541A9C5028A0BCDB14F851EC75971113D635FDEE0A93C85C3BE476FBCC1;
defparam sp_inst_18.INIT_RAM_34 = 256'h54F9318D0C53BBF084FA2725A842D0ACCD6C92633025E2B71DB975D28232EB7B;
defparam sp_inst_18.INIT_RAM_35 = 256'h8883FAF5068A5A7D64BE25BA89BA646E554732061B5102A8D80FDF2AC45DE119;
defparam sp_inst_18.INIT_RAM_36 = 256'h8D8768069C70B7E9F4AA889DA761B2466022259ED12BBC00FE5695B72401B82B;
defparam sp_inst_18.INIT_RAM_37 = 256'h79EAA00F3AF05E6FD5179E22E976B5B9D14742F042A1775A72E38D5EC6055506;
defparam sp_inst_18.INIT_RAM_38 = 256'hF3ACDA4D9DBEE7045B6C9E16553FFD37293A2339B00FFE9589DD48D81E99F0AA;
defparam sp_inst_18.INIT_RAM_39 = 256'h0E7C6A95555A89EC41551B4FDB8B5CFFAF010EAAC40EA619D414B301E0405F67;
defparam sp_inst_18.INIT_RAM_3A = 256'hF00FB3C0FD55287681A71E0BEF1CDC264A53301E269EAF60B32991509140EEB7;
defparam sp_inst_18.INIT_RAM_3B = 256'h5CF9916DAF33DEB9005593F1588BDAA40000055B8A2CF554B53086D7EE617498;
defparam sp_inst_18.INIT_RAM_3C = 256'h055AC5C47F10342E126DDF8AD5E9B28403FFCD6FEF009CB7786AD6D33698283A;
defparam sp_inst_18.INIT_RAM_3D = 256'h0EA90C2E7E6273B741DF607C9894BEEEB3CD647D79BA405503C056C669594000;
defparam sp_inst_18.INIT_RAM_3E = 256'h5084E5AA55690005AAAAFF2E50000556B5D70CB4CBFA9CD71753419E56D10EAD;
defparam sp_inst_18.INIT_RAM_3F = 256'h130F3812A3D058B42428FDD2A962FAA396E4EB95BC3ACA471C5D96DC1B2BB6FE;

SP sp_inst_19 (
    .DO({sp_inst_19_dout_w[29:0],sp_inst_19_dout[9:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9:8]})
);

defparam sp_inst_19.READ_MODE = 1'b0;
defparam sp_inst_19.WRITE_MODE = 2'b00;
defparam sp_inst_19.BIT_WIDTH = 2;
defparam sp_inst_19.BLK_SEL = 3'b010;
defparam sp_inst_19.RESET_MODE = "SYNC";
defparam sp_inst_19.INIT_RAM_00 = 256'h12AF001A1A0305AA96A93EA9A95555BC3001195500154000053E4290DABFF940;
defparam sp_inst_19.INIT_RAM_01 = 256'h555540055550F3F9014006AFFFFAA9556AA40040005550006FFF9000000056A5;
defparam sp_inst_19.INIT_RAM_02 = 256'h0000005554003FFF900005005A9550B575DD967C005556AA539AA51555AAAC00;
defparam sp_inst_19.INIT_RAM_03 = 256'h255105555AAA54AA95055AAAFF05555555040694FA640154C7FFEAFFFE555A90;
defparam sp_inst_19.INIT_RAM_04 = 256'h00150394057D2FDE4163AF8169000155555555002FFEA40014056A96D00AA952;
defparam sp_inst_19.INIT_RAM_05 = 256'h55001AFFA5155005A95BF5A91AA741A415AA55AA54FA55555AAF000555596950;
defparam sp_inst_19.INIT_RAM_06 = 256'h555A00FA555556AFC00F056AA45040C568A4047DFC92F39732D6A90155140551;
defparam sp_inst_19.INIT_RAM_07 = 256'h46A4F146AA9D97A6A940145400001550056A54155056A96FB993C56A315A56AA;
defparam sp_inst_19.INIT_RAM_08 = 256'h4000556AA96A9A96AB1BBBC656BA940554E9555556ABFC3EC15AA35140067F82;
defparam sp_inst_19.INIT_RAM_09 = 256'h5555556A3FF100CAA310411552826B90C7A6A969642AE400016A95A519554104;
defparam sp_inst_19.INIT_RAM_0A = 256'hA968945950555AAAAAA995555414500055AAA5566A694EA2F81556A9940514AA;
defparam sp_inst_19.INIT_RAM_0B = 256'h5565901AA4EA105056A4005403FA555555AAC00301F69F7A4000530283A462AA;
defparam sp_inst_19.INIT_RAM_0C = 256'hB24CC53D5056A500C54F30093BAF96F79055016AAAAAAAAAAAA5A5400055A6A5;
defparam sp_inst_19.INIT_RAM_0D = 256'h15AAEAA9AAAAAAA9A555556A5565156589A16F8A8145555553C543FA95565AAA;
defparam sp_inst_19.INIT_RAM_0E = 256'h8BE4041BF905A90043EA9696AAAAFC55154555315A406A40EDB4DE6A969E5040;
defparam sp_inst_19.INIT_RAM_0F = 256'h403FC6406AA4CB658ABAAA2900705AA955AA9516AAAA55555555156A555A9396;
defparam sp_inst_19.INIT_RAM_10 = 256'h95556AAA9500055515556955AA8E6DA9502AFD0016A43FFA955AAAAAB4066595;
defparam sp_inst_19.INIT_RAM_11 = 256'h6A40141A4FFAA55AAABFEC50464C0FFAC55605902F256C6543940175A954015A;
defparam sp_inst_19.INIT_RAM_12 = 256'hA52C55D61AAEA9000066A50000056AAA55AAA405554015406A4AC6F9EB14002A;
defparam sp_inst_19.INIT_RAM_13 = 256'hA56AA90001515A8A687F8F00C01A69002A0593EAA956AAFFCFD901ED13E60055;
defparam sp_inst_19.INIT_RAM_14 = 256'h193EAAA5AAFFF00655AF0E985693152AB0F211555500005695005401A96A51AA;
defparam sp_inst_19.INIT_RAM_15 = 256'h00000000005201400006F7C691AAA9A96A5A00556FE4AA8B950040C550057F90;
defparam sp_inst_19.INIT_RAM_16 = 256'h4D45AB9A4A9D550193C00003D9BD3D4FBFFD96BFC501192AE9546364BCBA575A;
defparam sp_inst_19.INIT_RAM_17 = 256'hEA6BF672103A665EFC7AA12E4A055500000000113C003F169ECBA6AAA5A5A57F;
defparam sp_inst_19.INIT_RAM_18 = 256'h000D0FF00006A5BFEAAAA56690BF81415506B9EA0FDBF80F03C2AB1BDE9CC260;
defparam sp_inst_19.INIT_RAM_19 = 256'h6E0E001E6D00C1BCFAADB3A04EC26FAAC01967AA269B54E97EC4D95054000000;
defparam sp_inst_19.INIT_RAM_1A = 256'h193AB9AB6498A74F640B54000001400850FF0002ABFFAAAAA455956A54069550;
defparam sp_inst_19.INIT_RAM_1B = 256'hFFF156A5005AA4155501506941511A40C5181900151AE2AB068503C4EAFA6143;
defparam sp_inst_19.INIT_RAM_1C = 256'h94030EAF6E2A450559143EABEB143C905A4EFB95AD7793FB55000000000B140F;
defparam sp_inst_19.INIT_RAM_1D = 256'h655675DC6C00554000000057F001B92B00000015A40000544195385405564159;
defparam sp_inst_19.INIT_RAM_1E = 256'h5555940440541A47DEB155692B0503BF5EA98B8A958F0008B3AAC2B653696DF2;
defparam sp_inst_19.INIT_RAM_1F = 256'h97B472443FC03AFEA17A29B8748D6AA96C2591C40000000000573FDFFF930000;
defparam sp_inst_19.INIT_RAM_20 = 256'h556200000000001283DFFFA640013C059014003069BFF8DB00102730F001F8EA;
defparam sp_inst_19.INIT_RAM_21 = 256'h0005A6FFEA9EAC003BED3C53FD8AB9D50C4670C0FFFFFB64B2936535BB3C1F50;
defparam sp_inst_19.INIT_RAM_22 = 256'h595450FFD7B69275956824169004959540154000005254EEEE6BF0003F168000;
defparam sp_inst_19.INIT_RAM_23 = 256'h5240000114E9557F8001056D000000066FFFFE8A69C53FF1C0E665D5D76B03C6;
defparam sp_inst_19.INIT_RAM_24 = 256'hE3FA83C00FD2FD89561EEEC031A9955655553C0F6A20A316905EF155A5A6AC5A;
defparam sp_inst_19.INIT_RAM_25 = 256'h3C50FD577B95E64D5B77AC3EFFFAE8E40001D5C53C6AC3004CF4064000696FFF;
defparam sp_inst_19.INIT_RAM_26 = 256'h9540E853B1401BCD6A554195BFFF0FEBBE4CC0FFE3DFA6671A3C194655A05555;
defparam sp_inst_19.INIT_RAM_27 = 256'h6C3FBEBF09A1270194F05A4FF15454000F1932A88A1605B95904FFEA503E4001;
defparam sp_inst_19.INIT_RAM_28 = 256'hB94669C24051959FFE403EFF500095443B40B0F17DC029A52A90FFF9FEA7FA4F;
defparam sp_inst_19.INIT_RAM_29 = 256'h842ED0065141694DC6FBF9EFFE3FABFFAB9575D98F074F03F62F3F15A40C6969;
defparam sp_inst_19.INIT_RAM_2A = 256'h5F0A00D80000338A93C155414C558A7C9A268057615E955A50FE900059444A10;
defparam sp_inst_19.INIT_RAM_2B = 256'h4414A7AA55AAA939500039A94F001BF9C02E85CA8F9568B794BFFB5A5556FFAE;
defparam sp_inst_19.INIT_RAM_2C = 256'h5A6AA7BEAAF9A3FFC9BE9D899BEA24E7FC67000303781A3F567E724168684693;
defparam sp_inst_19.INIT_RAM_2D = 256'h00030DB026319642050553F2812DD067EF56AAAA5A785000746BBAFFFF8C4005;
defparam sp_inst_19.INIT_RAM_2E = 256'hAAAAA94940007E410054EE54004D65A6FF8E56AA4FFE66954BD3A581B04FCC9D;
defparam sp_inst_19.INIT_RAM_2F = 256'hAAA5DFBD9A597F69660BFFFC0C73310330959D1965819064054F29558E466DD1;
defparam sp_inst_19.INIT_RAM_30 = 256'hA41AD643C5400FC1ADE3CAECF617AAAAA93914013E915E0188DB0000C55BAAF9;
defparam sp_inst_19.INIT_RAM_31 = 256'h140178FC2317F1F4010055ABBABE9EAF506DB99AF4EE5CA3CAEFFD85692E682A;
defparam sp_inst_19.INIT_RAM_32 = 256'hE54FDAE532CAFF0FF2703BFC5B8250F19A80C53CFAAC4F197D415975AAAAA4E5;
defparam sp_inst_19.INIT_RAM_33 = 256'h4313AAAAF1EEF8C6A0455AA55390140168054EDE3600000196BFBEAABDED4C17;
defparam sp_inst_19.INIT_RAM_34 = 256'h5F515E0C10065AAFBFAAEAE4013E563E3B91CA33340AAD3001AA90500043C57C;
defparam sp_inst_19.INIT_RAM_35 = 256'hA0D2C00551516AFFBF7140003230000EAAAAAF67068F642EC150F940150166A5;
defparam sp_inst_19.INIT_RAM_36 = 256'hA6B10F78ABFE5AAA550015015EA54BE4941A80286FEAABFFAAAA0129A8FBB05E;
defparam sp_inst_19.INIT_RAM_37 = 256'h3852AFFAEAAFFAAAE39A96A0EDB38EAFC40F5056532EDC8304F01500C03AAAAA;
defparam sp_inst_19.INIT_RAM_38 = 256'h430FCDAEA7850050270C0FEAAA956AAE0032DA97055000001501551265A6A52B;
defparam sp_inst_19.INIT_RAM_39 = 256'h0FF7000000001501570193298377AA19AAFFFAAABFFAAA796AAA040F363CE31C;
defparam sp_inst_19.INIT_RAM_3A = 256'hAFFAAEBFABE796955920DF57E5C241A854A6AE5C40018C4002AAAAAAAAAABC4E;
defparam sp_inst_19.INIT_RAM_3B = 256'h2E1100060030FAAAAAAAA95AABC0C00000000000154107AA55A9311AB4ABAFAB;
defparam sp_inst_19.INIT_RAM_3C = 256'h0000150142DAAE56614046BABDA2AEBFFEAABAAA75AA3377C1F4EA60005676E1;
defparam sp_inst_19.INIT_RAM_3D = 256'hFAAAA49509FCAA5D0EEB917D68859F0C05670000EAAAAAAAA96AAABF00000000;
defparam sp_inst_19.INIT_RAM_3E = 256'h0013AAAAAAAAAAAAAAAAFF0000000000050056A6AE60711969FAE0B46FAAFAAB;
defparam sp_inst_19.INIT_RAM_3F = 256'h55B287D1B068EFAF9BFE3DBEAAAFAAA9A57918F30F3A3E9EE91495527C405A30;

SP sp_inst_20 (
    .DO({sp_inst_20_dout_w[29:0],sp_inst_20_dout[11:10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11:10]})
);

defparam sp_inst_20.READ_MODE = 1'b0;
defparam sp_inst_20.WRITE_MODE = 2'b00;
defparam sp_inst_20.BIT_WIDTH = 2;
defparam sp_inst_20.BLK_SEL = 3'b010;
defparam sp_inst_20.RESET_MODE = "SYNC";
defparam sp_inst_20.INIT_RAM_00 = 256'hDC088020D7D6FDDD557FC0A28A0022ABEDF5FFD7DFDFD55F5DC88A889DDDDF5F;
defparam sp_inst_20.INIT_RAM_01 = 256'hFF7D777DF5778E80A02057FFFFDD7FDDD7DDF5D555DD77DDF7FDDFFD7D75D5F7;
defparam sp_inst_20.INIT_RAM_02 = 256'hFFD55DD7F77FFFF75557DFDFFFDDF52D4892BFE1F5DFDFD7F600820028A029DF;
defparam sp_inst_20.INIT_RAM_03 = 256'h5DD75DF5DDDFD5A00220000820D577DDD7DDD75F82A808AA1FFF5DFDD7577F5F;
defparam sp_inst_20.INIT_RAM_04 = 256'h75D5DC0A0AA27FD2888FF5D55DFD5FFF777775777FFFDF5F7FDF57FD777DF75C;
defparam sp_inst_20.INIT_RAM_05 = 256'hDDFD7D55DF7D5775DDDDF5DD555677DF57FD7DDDFF2AAA000022DFDD5FF7D55F;
defparam sp_inst_20.INIT_RAM_06 = 256'hD7FDDD020280000A3DF8DF5757F5F537F7AA2A227D8A8C2A4DFF5DF5DD5FF7FD;
defparam sp_inst_20.INIT_RAM_07 = 256'h8882DEB5D77A00FF77FDDF5DDFD5F7D777FDDF7555757F7FFD76BFF74DD7DDF5;
defparam sp_inst_20.INIT_RAM_08 = 256'h5F75F777DDDFF5FE207FFE15D5FD57FD772008A80000896815DFFE5DFD5DFE9C;
defparam sp_inst_20.INIT_RAM_09 = 256'h008000026AAFF5B774FFD7F5DE34A2205ADF77FFA25F5FD7FF7D7F7F7DFDD7FF;
defparam sp_inst_20.INIT_RAM_0A = 256'hFF75289F5F5F5DFDFDD777D7DDF5F755F5FDD5DD77D7D00FFDF5FD7D5575D580;
defparam sp_inst_20.INIT_RAM_0B = 256'h557F5FDDDF0AF55557557D7FDE00000000081FD4F5077255F575FE569C804FDD;
defparam sp_inst_20.INIT_RAM_0C = 256'h8FF13FC15D7D57579DDAE7F2EF7DDD5400977FDDFFD55F55FD775F775D5D7755;
defparam sp_inst_20.INIT_RAM_0D = 256'hD7DDD575DDFF7F777DD775F7D77577FFD88DFFD09DFDDD7F5435FEAA82000008;
defparam sp_inst_20.INIT_RAM_0E = 256'h1FFD5F7577D75F75FEAA02000002815D5FD77FC75F57FFD58BC83575FDD20A1D;
defparam sp_inst_20.INIT_RAM_0F = 256'hDD4A3777D5F715E2157FFD420825FDFD55757FF55FDF5FFFF7FFFFDFFD7756AA;
defparam sp_inst_20.INIT_RAM_10 = 256'h7D5FF7FF55D7F5D5FD5DF5FD5DF883577577FFDF7777680080000002ADFD577D;
defparam sp_inst_20.INIT_RAM_11 = 256'hFF7D75F7D222000200282BDF75D1F2023FD7D75DFFCA2B7FD62A02275775775D;
defparam sp_inst_20.INIT_RAM_12 = 256'hF54BDDA8A80000A808A57D5DD777D75F7D5DF5D75FF5777DD558BD5580575557;
defparam sp_inst_20.INIT_RAM_13 = 256'hDF75D77F7D7D5FF009DF50F7B75FF77FD5FD74882200000A921D57A976A0F5DF;
defparam sp_inst_20.INIT_RAM_14 = 256'hD56020000000257D57A0D023DFDEF7CA07A520A8A088280DD5DDDDF7FFF5DDFD;
defparam sp_inst_20.INIT_RAM_15 = 256'h828280222A8FD57DDF5DF635F5FD7F755D755FF757DD803F75D5F71D755DDF77;
defparam sp_inst_20.INIT_RAM_16 = 256'h5155DFFF70A1D5FF5635D77C37F7E158A0AA0028157FFFE02AA976D501C288F5;
defparam sp_inst_20.INIT_RAM_17 = 256'hA0028DEFF5EA0A0A09E22F417AD580200000028F63F5C87FFABDDD575D57D5DF;
defparam sp_inst_20.INIT_RAM_18 = 256'hA209D205F75F57FF577755D7D77FFD75DD7DFF08FA3DD7F2DC16287DD2951607;
defparam sp_inst_20.INIT_RAM_19 = 256'h55F85FFF7D5F3757882BD6D7D8B62000BD75748060285FA20A979DFF0A0200AA;
defparam sp_inst_20.INIT_RAM_1A = 256'hD74A8002F7880AFA7FFAA28200A02203FD82F577D7FD7F775555FFD7D55F57FF;
defparam sp_inst_20.INIT_RAM_1B = 256'h8227FF57FF75557F5F77DD75F77F5777377FDD5FDD7F7622DFFFDC9D808A0F56;
defparam sp_inst_20.INIT_RAM_1C = 256'hD75ED022DFE01FF57DF5C002A875C9DDD000288829EFF4020202002820207778;
defparam sp_inst_20.INIT_RAM_1D = 256'hA02807BF2BF7A0A0000008828755DDC0FF55D557F7F75D5F7D576155DF7FD57F;
defparam sp_inst_20.INIT_RAM_1E = 256'hD77D7D555777DF75F285775D6077DCA258A897D817D0D552A40036A5DEF74B04;
defparam sp_inst_20.INIT_RAM_1F = 256'hAADFEDFF68BDC000ADC2FF5747102282A3DE0A17022000000AAAC217FFD6755D;
defparam sp_inst_20.INIT_RAM_20 = 256'hA22E8A00A00008A0D61FD5DCDD77E17DDDFF7FEDD7FD5F00D7FDE0E587DDDF02;
defparam sp_inst_20.INIT_RAM_21 = 256'h557FFF7DF7D023F7E289C3F6ABD8229D73DF6F178000A8D70F5ED7400A6372D5;
defparam sp_inst_20.INIT_RAM_22 = 256'h57DFD5803E257DE57D575FDDDDD782892A8888000800D71D775687F54AFDFD7F;
defparam sp_inst_20.INIT_RAM_23 = 256'hD6AAA8A8DDB7D7F63577757DD75FF5DFF5FF775A0A17EA0D178A2217287CD4B7;
defparam sp_inst_20.INIT_RAM_24 = 256'hF4081E17DABE03D20AA949FD65577F5D7DFF61DA7FC55C77FDF885D708A889D5;
defparam sp_inst_20.INIT_RAM_25 = 256'h4B7D0954AD7787DA82DC8142FFDDDD8222AA1715E9DE347D5155D7F7F5D7DFD7;
defparam sp_inst_20.INIT_RAM_26 = 256'h3777815EA5557D73D5F7FF7F7FFD50AAFD539F8027D88AAADDE1D7DFFFD57D7D;
defparam sp_inst_20.INIT_RAM_27 = 256'h09C22A00582ADE775FAFFDF807DDF5777AD545773F560A8A9D77FFFD7740A00A;
defparam sp_inst_20.INIT_RAM_28 = 256'h77FF751608A097F2FFF5422A28283D7D62F72525F59575FD75775FF78AA5F572;
defparam sp_inst_20.INIT_RAM_29 = 256'h15FD7D7F57D57FD815FE02BFDF6880A028A88529FAD55254276A487FDDF1D5FD;
defparam sp_inst_20.INIT_RAM_2A = 256'h897F5F9FDDF74C17761DF5FD5B57976375E02A0A057AD5F577288828377DF0FF;
defparam sp_inst_20.INIT_RAM_2B = 256'h8A230EBCFD777D62080827F7F2D7DF7F1DD5F5B5D28001FC837FF68A00A20A8A;
defparam sp_inst_20.INIT_RAM_2C = 256'h5FFF5E880A8AA5D7D8022B58A820433C21F4DFF45E7DDDC25563C77DCBF5F75E;
defparam sp_inst_20.INIT_RAM_2D = 256'h7D7C79402FE7F557F77FF405DDD7A028087ADFF75D62A8088F57FDFDF7715DFD;
defparam sp_inst_20.INIT_RAM_2E = 256'h5F77F7D88A0205F577D51DFFDD5BF55F7F78000037F7E2A01F5EA014877899D3;
defparam sp_inst_20.INIT_RAM_2F = 256'h80021F752882F76288528A8153E447FC4DDA9D7F7777FD5DDF50F5D7D00AC1A7;
defparam sp_inst_20.INIT_RAM_30 = 256'h5FD7F5DEBD77DA1709DC3D292FF45557DFC80200A7F552F737947555BF7555F5;
defparam sp_inst_20.INIT_RAM_31 = 256'h0A00AF89567D875F5755F5F5757F7820757D20AB5D82AB8C980801F7557FFD7F;
defparam sp_inst_20.INIT_RAM_32 = 256'h80BF5A2A8C982A72A5674229575775257FD71563A2015A7F6BF75555F57F7F80;
defparam sp_inst_20.INIT_RAM_33 = 256'hFCDCA020872B7FBD5DF3DD75F6A88008A7D778BD6DFDD57DFF7F7DD7F5217B74;
defparam sp_inst_20.INIT_RAM_34 = 256'hD0DDDDD3FDFF77FFFF5FD5FF554002FF4A8A12CEC5FA09C5FFFFFFFFFD74374B;
defparam sp_inst_20.INIT_RAM_35 = 256'h279697D57FFD7DD7FC8F5F5D6DCF7D52A028A856FDF057633DD7080A8A08A5F5;
defparam sp_inst_20.INIT_RAM_36 = 256'h8AA5F87F082D82A0202AA08A81FD757775DDDF5F7FDDD7FF5F557DE001FD6D02;
defparam sp_inst_20.INIT_RAM_37 = 256'hFD7D5FFFDF5FD57FDC8A822FD8AE92A2B7705777DC5DFFB6DD855DDDB5420A28;
defparam sp_inst_20.INIT_RAM_38 = 256'h54D8129DDE955DFD54F35A02A222A2AA7DCF5756220A02802200A155F77705DC;
defparam sp_inst_20.INIT_RAM_39 = 256'h5888A0A000002882A0FFF4571ED6D5777FDFF7FFDFFD77C80202D8F84DC30671;
defparam sp_inst_20.INIT_RAM_3A = 256'h5FF5F775F7FE02008B67357EA2B7FF7D7FA558DB5577537FDC20288802A82B50;
defparam sp_inst_20.INIT_RAM_3B = 256'h5875F7FF7D670A22A00AA2A0AA3797DD0000000228A0205F555D6DDD57DF75FF;
defparam sp_inst_20.INIT_RAM_3C = 256'h00020880A057557F67755557D587FF5577FFF575C2008C0E375D82277DFFED05;
defparam sp_inst_20.INIT_RAM_3D = 256'hF7FD5D20DA0380F21780DF437F3F58717FD475F72A28800A0AA0A828FDDF0000;
defparam sp_inst_20.INIT_RAM_3E = 256'hDFFE0A0002AAA000AA0002D580000000A88200D57ADDCF7FD7FD55D7DD77FD7D;
defparam sp_inst_20.INIT_RAM_3F = 256'h025777F545F73FF777D5E1FFFF7757FD55E9632EF8E27D7A1DFFDDDDC957554D;

SP sp_inst_21 (
    .DO({sp_inst_21_dout_w[29:0],sp_inst_21_dout[13:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13:12]})
);

defparam sp_inst_21.READ_MODE = 1'b0;
defparam sp_inst_21.WRITE_MODE = 2'b00;
defparam sp_inst_21.BIT_WIDTH = 2;
defparam sp_inst_21.BLK_SEL = 3'b010;
defparam sp_inst_21.RESET_MODE = "SYNC";
defparam sp_inst_21.INIT_RAM_00 = 256'h98001021EFFD6310420D90FDA400606A42A26903AA84FFC0189E9421C27EF773;
defparam sp_inst_21.INIT_RAM_01 = 256'h03EA99750697B00B06956447BFE33E0070EE950055198BBCBFFF8F56FC06B7E7;
defparam sp_inst_21.INIT_RAM_02 = 256'h0000550B9CEADFFFD594BFC1B7E0EEB1FBEE6608C865B7173DEAA4001BFEAD6B;
defparam sp_inst_21.INIT_RAM_03 = 256'h95401800C41357DAA9400550F3DC3EBFC270B6F9540D02A9EAFFE6FFBC436F87;
defparam sp_inst_21.INIT_RAM_04 = 256'h9BDA007405AFCFC2FBD51FC2F9905555AE4B9229DFFAEAE5FFC66FEB0E6A17F1;
defparam sp_inst_21.INIT_RAM_05 = 256'h137A56AA9A31031CCF87A86475B0CDAB61AA82D303791BE4000567DBFADAB8FA;
defparam sp_inst_21.INIT_RAM_06 = 256'hDF2F00881FE4000600FF6B759BE695654A9C04B2FFBE146D71A308406AA56E46;
defparam sp_inst_21.INIT_RAM_07 = 256'h4410B703A5808A0B3B4F6AFA6A55C493116C5D0B55B60D8BB2913B19BDA8C469;
defparam sp_inst_21.INIT_RAM_08 = 256'h53F65A1FC945D594A276B1DAB2FF6D7647641B900006FC3A1C4BE1E29577BDA4;
defparam sp_inst_21.INIT_RAM_09 = 256'h000000003FEC350B908FEABA35935DDDD35D1728D8CC71031B55554EC5E50BF0;
defparam sp_inst_21.INIT_RAM_0A = 256'h54173A90206C710150C3E9060903A9B1F6FFB96BC7D96FCFA91B6DAA93F17A90;
defparam sp_inst_21.INIT_RAM_0B = 256'h15AA2EE284DF5D50CB0E9753C8E400000001D412F61A698F2A5A505FE96CD651;
defparam sp_inst_21.INIT_RAM_0C = 256'h7911CC844DE7279488C4EC94066F8DF0397E41D8C5555000FF9AE2940C6C5AF9;
defparam sp_inst_21.INIT_RAM_0D = 256'hDC81C5450FAC003EE500401A15A9F06AF9745B51D504C006496137A400000001;
defparam sp_inst_21.INIT_RAM_0E = 256'h43D1C32F9F0BA4EFE4E500000000C61380000B81FE24D9DEDB34EE19827CE455;
defparam sp_inst_21.INIT_RAM_0F = 256'h014FD0CF6A4B968401AA95A355758BF9C6F1240B155E90015400BF2AC1AF6DD6;
defparam sp_inst_21.INIT_RAM_10 = 256'hE6AAF0539E5AFFAABFC11A9655C4255A3A6FF92BCAE7413A000000000CA2BF25;
defparam sp_inst_21.INIT_RAM_11 = 256'h6568C51F37E940000001DA509DCC03348BEBF1755E368900E779196BC278F618;
defparam sp_inst_21.INIT_RAM_12 = 256'h431473453C5A93541513489FC55DC5A4D210DD2F5395F3EB2FB089F727DCAA7F;
defparam sp_inst_21.INIT_RAM_13 = 256'h32DFBD2AEBEB7102B3AFFF125AFCFAE2F44621E5400000007E5F704FBB82B1A6;
defparam sp_inst_21.INIT_RAM_14 = 256'h7DB90690000012F4D7FDC121823E1ECA3947165FAE1505509E0C15F9696F0780;
defparam sp_inst_21.INIT_RAM_15 = 256'h014400040553903CC0CCFA7B82804873C0ECD1AC8BD2563EF23A6438E78E5FB7;
defparam sp_inst_21.INIT_RAM_16 = 256'hBE69867C334158939E065B190F7CFEC45F4000508D2B9E2B1B52B38DB9EA66BB;
defparam sp_inst_21.INIT_RAM_17 = 256'h40008F54C57A1FA2B9B71E3680DBFF800000011786F0E04BC2E788A459E0F9AF;
defparam sp_inst_21.INIT_RAM_18 = 256'h0003395BFD6DE5BFD04D5866E03FC0E4BF49A026AD9EF640BF3EB2236877EB69;
defparam sp_inst_21.INIT_RAM_19 = 256'hECDE241FFED2CBF9514922C7AEE005004B142B6A5A9FC882E447AE76FA400000;
defparam sp_inst_21.INIT_RAM_1A = 256'h093A6C70103DF58A0FEDA9000005400DA2000E4F6FF996035B16A599E1D23FE5;
defparam sp_inst_21.INIT_RAM_1B = 256'hCE87C6E26D265A55BEA0F5ED405B74B92399D4E68566B140D7C1F463B0241474;
defparam sp_inst_21.INIT_RAM_1C = 256'hE0C9A40BE80C19DCA949CC05D3CDFFA6FD0F3AD6FB6A3BF7A9400001014857D1;
defparam sp_inst_21.INIT_RAM_1D = 256'h5E4B996DCDAB5A4000000157AA18D2A01B39B0763354A6C0E0E5CD2A6BD00115;
defparam sp_inst_21.INIT_RAM_1E = 256'hCD32160040AE528A919D5AF4F855742F97CEC740786C667336008642A007D456;
defparam sp_inst_21.INIT_RAM_1F = 256'hEA2BC5E3E64EB01010CA59354F0C22BEBB0978E255400000005325C7FF6A4001;
defparam sp_inst_21.INIT_RAM_20 = 256'hFFCC505500000053D2EFFFA7E00B54E3BD050007E9DBE168855D12E42A3DFF7B;
defparam sp_inst_21.INIT_RAM_21 = 256'h5AA20CFBEA66B84E914CF8223E0FC3BEE8B44123400594DC8F996261B087D951;
defparam sp_inst_21.INIT_RAM_22 = 256'h1FCE537032831E0ED3ECC9847658D0F0D06B500000923C3FD976A41C56D6055A;
defparam sp_inst_21.INIT_RAM_23 = 256'hF5800101894D84D52E5A7F62F801EA9027FFFD391005C9B4DAB16A021587BFD7;
defparam sp_inst_21.INIT_RAM_24 = 256'hD685FDBE073CC9CDA415D030327E3AE7FF74D20AA0B2FB88CB098BBD40CD22C5;
defparam sp_inst_21.INIT_RAM_25 = 256'hB13BC096ADC3073BC8EE07E8BFFAA2DD40000D0B97C614069BB77DA96CFD4BFE;
defparam sp_inst_21.INIT_RAM_26 = 256'h6AAEE72C190006C971DD5125BFFF89D93D6583B042FB0265BD7E84F2CED75BEB;
defparam sp_inst_21.INIT_RAM_27 = 256'hB43A7D8311E17F019DF1AAC424819A0B9BED903AEF2DAC86D407FF9639484000;
defparam sp_inst_21.INIT_RAM_28 = 256'hBE8E6185EABB24C0F8954EFED001BA9A7624180EA6AA907F3CD2BEA6A277F9F4;
defparam sp_inst_21.INIT_RAM_29 = 256'h3466B91A00D4F89874F348EFF8BA6C15478F0E53AA1FDEF9AD5AAB7819482482;
defparam sp_inst_21.INIT_RAM_2A = 256'hF30B3E8ABF9406B3730AC2616206AB515FFCC5CF51550FC5383AE001482A710E;
defparam sp_inst_21.INIT_RAM_2B = 256'h05B295FAFC5454B7E0012DA8A0C3317304350367FB400FDA463E53F001466929;
defparam sp_inst_21.INIT_RAM_2C = 256'hAD80AEF401C809FF93D6420E4945C0EE98E2FAA4076BEA82C4D24EF7A53F24C9;
defparam sp_inst_21.INIT_RAM_2D = 256'hABE50766871BB54687AF67CC71E600206FE6155415C69001477FCC05FEC0003E;
defparam sp_inst_21.INIT_RAM_2E = 256'h554554D75005323BE5A93F461001390FAF8800001BFC8B8077FD40FEA0554878;
defparam sp_inst_21.INIT_RAM_2F = 256'hE000256CAB097D98F7EB540029439DE90491C07CD79D9F6C76907217B70E4AA0;
defparam sp_inst_21.INIT_RAM_30 = 256'h3FAB1D59DCBF0F1BF63D7E65F02E55551373A4062A76E8C20FDF0000970BFFF8;
defparam sp_inst_21.INIT_RAM_31 = 256'hA4061E380570435A000AC86FFFFE910BAB9B2DDCF858E3FB11401DB22D22115F;
defparam sp_inst_21.INIT_RAM_32 = 256'h643FC88A2A769449675841ADADB892521C59B0DB3EC6E0DA056D593E05404DDE;
defparam sp_inst_21.INIT_RAM_33 = 256'h3443F03FCB52FC535B02C140E62569023A5A9DCC92784063ADFFFFBEBF5E38C6;
defparam sp_inst_21.INIT_RAM_34 = 256'hBF6E36D7C97CCBFFBFFAFFBCF27E01EDFA20BBE4F6506DD5C7BFEF6A97399632;
defparam sp_inst_21.INIT_RAM_35 = 256'h2E9A4EAFF977863EEA55FB0FDA6AFAD70541C1DF249C884A06A9349069026253;
defparam sp_inst_21.INIT_RAM_36 = 256'h4FF764E6F15DC5553E406E01536CE57841FA04616FFBBFFFBFE4975015138467;
defparam sp_inst_21.INIT_RAM_37 = 256'hB3A6FFFFFAFFBFFFCD4002BCDAE9C7071D4C0B9C0A6FDD8C80AC23FFA1405541;
defparam sp_inst_21.INIT_RAM_38 = 256'h7AF365CEEC594C0F63ABFC550543D8C369FB1B935AA554006E4144CE953BD1AD;
defparam sp_inst_21.INIT_RAM_39 = 256'hA513050000006F4095A83EF109E0588DEABFFEAABFFFE9581469C0A11320D883;
defparam sp_inst_21.INIT_RAM_3A = 256'hFFFFFEAFFFDA404004FC0A94D0E21FA64410CC6D8FE2F028801941504001C091;
defparam sp_inst_21.INIT_RAM_3B = 256'h9C1CAB123F9C9054555003F0005A1415000000006F4099EA15C8B6DB2D7BAE5B;
defparam sp_inst_21.INIT_RAM_3C = 256'h00006B41806DC606614BD7BFBA03FFFEAFFFFEAF3800200246F82A510B62BC92;
defparam sp_inst_21.INIT_RAM_3D = 256'hFEAA9F848CFFD2FA37BD8184699ED34C0713FE84405555500FF0000150C00000;
defparam sp_inst_21.INIT_RAM_3E = 256'hBA2700555400F000000053C0000000001B409B16788F596559F7C02C37EFFFEB;
defparam sp_inst_21.INIT_RAM_3F = 256'hA6271D5EDB154FAE217C457FFE9AFEA5F02CCEE41F33AE548F72269E13EA1C14;

SP sp_inst_22 (
    .DO({sp_inst_22_dout_w[29:0],sp_inst_22_dout[15:14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:14]})
);

defparam sp_inst_22.READ_MODE = 1'b0;
defparam sp_inst_22.WRITE_MODE = 2'b00;
defparam sp_inst_22.BIT_WIDTH = 2;
defparam sp_inst_22.BLK_SEL = 3'b010;
defparam sp_inst_22.RESET_MODE = "SYNC";
defparam sp_inst_22.INIT_RAM_00 = 256'h655500056A545AFFAAFA550000000555555AAAA9556A556AABA501402FFFFE94;
defparam sp_inst_22.INIT_RAM_01 = 256'hA955555AAAA95AA400005BFFFFFEEAAAAFA555555556A4016FFFF40001555AA9;
defparam sp_inst_22.INIT_RAM_02 = 256'h55555555A5007FFFF90000155AAA550A90646A9116AA5AFE9500000000000155;
defparam sp_inst_22.INIT_RAM_03 = 256'hBAA556AA6BFEA9000000000004169555695A5AAA555000001BFFFFFFFFA9AAA4;
defparam sp_inst_22.INIT_RAM_04 = 256'h556AAA4000147FF9001BFFAAAA5555555555A9407FFFF9000015AAAAE55AFEA9;
defparam sp_inst_22.INIT_RAM_05 = 256'hA9406FFFF9455456BABFFAAAAFFEA6A45AAAAABEA940000000005415556AAA55;
defparam sp_inst_22.INIT_RAM_06 = 256'hA5AAAA5000000000550055AFF955555ABE500018FE41AA419BEAFA5555555555;
defparam sp_inst_22.INIT_RAM_07 = 256'h0154F86FFFF951FAE950555555556A545AABA555555AFABFFEA95AFF96AA6BFF;
defparam sp_inst_22.INIT_RAM_08 = 256'h540555AABABFFFA905AFFD6AAFFFE55AA94000000000014056BFF955555ABE69;
defparam sp_inst_22.INIT_RAM_09 = 256'h000000004001456FF965555AA9680150E5FBFEFF107BE95455AAAAA56A55555A;
defparam sp_inst_22.INIT_RAM_0A = 256'hFFFE402A9556AFFFFFBEAAAAA55400055AAAAAAABEBF9016F955ABFFA95AA900;
defparam sp_inst_22.INIT_RAM_0B = 256'hAAAAE56FFA50A5556AFA55A96500000000001554055BE5BA9555AAA415509BFF;
defparam sp_inst_22.INIT_RAM_0C = 256'h06951656A6AAE9556BA556A4AFFFFBFE4015556BBFFFFFFFAAAAA9555156AAAA;
defparam sp_inst_22.INIT_RAM_0D = 256'h16BFBFFFFAABFFEAAAAAAAAAAAAA5AAA9006FFE415566AAAA55A940000000000;
defparam sp_inst_22.INIT_RAM_0E = 256'h6FF9145BF955AA5555000000000015A96AAAAAAAAA95BFA556D06FFFFFE50015;
defparam sp_inst_22.INIT_RAM_0F = 256'hAAA56FA5FFF96F906FFFFF9400056AAA6AAFEAAAFFFAAAAAAAAA55AA6AAAE500;
defparam sp_inst_22.INIT_RAM_10 = 256'hAAAAAFFEA5555555556AAAAAFFA506F9406FFE406AA9554000000000165AAAEA;
defparam sp_inst_22.INIT_RAM_11 = 256'hFE416AAA94000000000001AAABA6A9956AAAAFEABF8016FFA9400005BE9505AB;
defparam sp_inst_22.INIT_RAM_12 = 256'hFE96AE4101555400000AFA501556BFFFAAFFA555A9555955AA956BFE4065006F;
defparam sp_inst_22.INIT_RAM_13 = 256'hE96AAA955555AFE405BF9054001BA9056FAAE90000000000006A9A56A9555AAA;
defparam sp_inst_22.INIT_RAM_14 = 256'hAA4000000000055BA906B9466AE5AA505A5B00000000000BA5515506FFFFE5BF;
defparam sp_inst_22.INIT_RAM_15 = 256'h00000000000A55411517FEAFE5BFFAAEBFAB5556BFF9005BE94040065416BFE9;
defparam sp_inst_22.INIT_RAM_16 = 256'hD006BFEBD406A505A40000556AFF56A51554000016956A959401A9BA569001AF;
defparam sp_inst_22.INIT_RAM_17 = 256'h000016966A95500456945686A56A0000000000050005001BF96FFBFFFAAAAABF;
defparam sp_inst_22.INIT_RAM_18 = 256'h000540000007FFFFFFFAFAAAAAFFE506AAABFE40501BFD00005405AFE56D1405;
defparam sp_inst_22.INIT_RAM_19 = 256'hBF50556FFE0015BE5556F9B95019000015AAA9559001BA5415696A9500000000;
defparam sp_inst_22.INIT_RAM_1A = 256'h6A955006FE4001A5F95100000000000154005001FFFFAAFEF9AAAABFA91AEAAA;
defparam sp_inst_22.INIT_RAM_1B = 256'h10006AA901AFF955555A556AAAAAAF95596FBE006AAFE9556AAA556E40000695;
defparam sp_inst_22.INIT_RAM_1C = 256'hA9105555BF916A56AABFA000006501AAA0059500069BE9550000000000015400;
defparam sp_inst_22.INIT_RAM_1D = 256'h50001A6E16AA0000000000000056BE400040055AE800001506AA51AAAAAAAAAF;
defparam sp_inst_22.INIT_RAM_1E = 256'h6545E40000001AABE416AAAA415A4000A4102FE56A9195A89400141A55BE9659;
defparam sp_inst_22.INIT_RAM_1F = 256'h01F956594065400006506AFEE965540005B8416E000000000000402FFFE40000;
defparam sp_inst_22.INIT_RAM_20 = 256'h0015000000000000542FFFF800005505900000006ABFFE416AA540064056F940;
defparam sp_inst_22.INIT_RAM_21 = 256'h0005FBFFFFE406A5000241A996E0146A015B40540000016516FAFE95555565AA;
defparam sp_inst_22.INIT_RAM_22 = 256'hAABAA940041AAB9BA96A796BEAAA0007000000000000956FFFFD0001001B9000;
defparam sp_inst_22.INIT_RAM_23 = 256'hA9000000657FBFBD0000406E0000001BAFFFFFD0006A5006154000BE41B8001A;
defparam sp_inst_22.INIT_RAM_24 = 256'hF9501555A45516A00107D7D545AAEAAAAA9500506F4AA46BA5A56AAA50115ABF;
defparam sp_inst_22.INIT_RAM_25 = 256'h404016A91BA95A9416B95555FFFFFE500000656AAAB8000001F80640016ABFFF;
defparam sp_inst_22.INIT_RAM_26 = 256'h1555559000001BE01FA506EAFFFFA501FF95695A5BE55001AA406A5ABAA4AAAA;
defparam sp_inst_22.INIT_RAM_27 = 256'h06955569A400A455A505AA5006BFA400506A5BE91AA901642AA9FFFFEAA50000;
defparam sp_inst_22.INIT_RAM_28 = 256'hAAA6AE6900006AA5FFAAA5550000155540400001BD002FE55BA9FFFE540BFF95;
defparam sp_inst_22.INIT_RAM_29 = 256'h056FD006AA56AA505BFD502FFF95015555506A46905650000640005BF901AABE;
defparam sp_inst_22.INIT_RAM_2A = 256'h0BAA40290000001EE801BE4695AA1A95AA4100115AA4FABFEA9500002A954050;
defparam sp_inst_22.INIT_RAM_2B = 256'h00065928ABFFFF9400001AAA5569AFE9001FE90AE40001B901FFFD0500005555;
defparam sp_inst_22.INIT_RAM_2C = 256'hAA6FF900001007FFE41406E0015556640168000000BEBE00BF46564641A99BA5;
defparam sp_inst_22.INIT_RAM_2D = 256'h000001E52E46AF96190654179A6E405695A0FFFFFFA4000019AABBFFFF900006;
defparam sp_inst_22.INIT_RAM_2E = 256'hFFFFFFA400000E9555551AA40001AAFBFFE000001FFF90001FE500141A901191;
defparam sp_inst_22.INIT_RAM_2F = 256'h00006FFF4000BF95005000000194010001BA7E5BBE91A5A50555AEA99401964A;
defparam sp_inst_22.INIT_RAM_30 = 256'hE41AEB901640505506E55A465FA9FFFFFE9400001E955015192900001AFFFFFF;
defparam sp_inst_22.INIT_RAM_31 = 256'h00001941645B55F400006BFFFFFFE40055BE5003FA55050450000299AAAEA96A;
defparam sp_inst_22.INIT_RAM_32 = 256'h401FF5501450555006955556AB815405AB9005004015556A9696FFFAFFFFFA50;
defparam sp_inst_22.INIT_RAM_33 = 256'h401405401546AA5AFAE6BFFFA94000000955502B9A400005ABFFFFFFFE414169;
defparam sp_inst_22.INIT_RAM_34 = 256'h50A6AE001007BFFFFFFFFFE50540007F954050555950025515AAA59000401A80;
defparam sp_inst_22.INIT_RAM_35 = 256'h4564655556956AFFBD15005006400014555515645B91BA96AAAA950000000AA9;
defparam sp_inst_22.INIT_RAM_36 = 256'h50055569055A15554000000006A65BEAA91BE56EFFFFFFFFFFFF554001FFEA04;
defparam sp_inst_22.INIT_RAM_37 = 256'hBDABFFFFFFFFFFFFF5000006F41524545551A5A6A5BFFE101501590005555555;
defparam sp_inst_22.INIT_RAM_38 = 256'h9554543FF915515068000155555415145506EAA800000000000002666AEA057E;
defparam sp_inst_22.INIT_RAM_39 = 256'h55500000000000000156956E507EFFBFFFFFFFFFFFFFFF90000060559A950565;
defparam sp_inst_22.INIT_RAM_3A = 256'hFFFFFFFFFFF9000002466FA9001A95A9550BB051500595411555555555551555;
defparam sp_inst_22.INIT_RAM_3B = 256'h6051005A40015555555554055555555500000000000001AAAABA451BFAFFFFFF;
defparam sp_inst_22.INIT_RAM_3C = 256'h0000000001EABEAA8555AFFFFE5AFFFFFFFFFFFFD00019196AFA4005505A4605;
defparam sp_inst_22.INIT_RAM_3D = 256'hFFFFF900600115A41E41A556A915A45155A80015555555555005555555150000;
defparam sp_inst_22.INIT_RAM_3E = 256'h00545555555505555555541500000000000000FAE5B5955ABFFFFAFAAFFFFFFF;
defparam sp_inst_22.INIT_RAM_3F = 256'h00FAEBE695A97FFFEFFF56FFFFFFFFFFFFD24105A594BFE57959EAA69555AB95;

SP sp_inst_23 (
    .DO({sp_inst_23_dout_w[23:0],sp_inst_23_dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_23.READ_MODE = 1'b0;
defparam sp_inst_23.WRITE_MODE = 2'b00;
defparam sp_inst_23.BIT_WIDTH = 8;
defparam sp_inst_23.BLK_SEL = 3'b001;
defparam sp_inst_23.RESET_MODE = "SYNC";
defparam sp_inst_23.INIT_RAM_00 = 256'hACCC2C8C0C6C6B6B8161200000010000002141616160606081C24485034040A1;
defparam sp_inst_23.INIT_RAM_01 = 256'hACAD8D8C6C6B6B8B8B8B6B6B8C8C8C8C4B4B4B4B6B6B6C8C8CAC8C8C8C8C8C8C;
defparam sp_inst_23.INIT_RAM_02 = 256'h182B2EB371B77A77B37235B6F3D234F3B8D9987BDC96708C29094BEEF00EEB4A;
defparam sp_inst_23.INIT_RAM_03 = 256'hA856766EEE70B137B85B78130FCA88CDB9BABB1D1D56F010731510AE91D75A36;
defparam sp_inst_23.INIT_RAM_04 = 256'hF775335292F2B477199756B75978D5129696B6B69676553515B7D6902FF877CA;
defparam sp_inst_23.INIT_RAM_05 = 256'h55B316D1AC1154942F2AEDD157D10C4C4914D7F8F7397A7336FDFEBEFF7CB97B;
defparam sp_inst_23.INIT_RAM_06 = 256'hA261400021210000002141616160606060A224A644814081E486206DBA78B4D7;
defparam sp_inst_23.INIT_RAM_07 = 256'hACAC8C8C8C8CACAD8C8C6C6B6B6C8C8C4B6B6C6C6D6D6D4D4C6DCD0D4C8BCAEA;
defparam sp_inst_23.INIT_RAM_08 = 256'h71B22F6C2B6CEE2FD35A11CC7598720C098C303230EC6BACADADCEAD8C6B6B8B;
defparam sp_inst_23.INIT_RAM_09 = 256'hD93BB9F633CDCA4B0ACA3136F1ACAF5535D06E55B7F12FEE953BF56E5592092E;
defparam sp_inst_23.INIT_RAM_0A = 256'h97F818D755149517B6B6B7B6967696D776357537F6F0ECB0F70B8A1398D8F9FA;
defparam sp_inst_23.INIT_RAM_0B = 256'h6B2D16F63289280F497A7AD77A35D478FF9DFFFF5C7C7CF59B5E9E9852CE2F90;
defparam sp_inst_23.INIT_RAM_0C = 256'h0021416161404040608123A685C24040A203E314BA78D5D45054F5125679128F;
defparam sp_inst_23.INIT_RAM_0D = 256'hAC8C8C6B6B6B6C8C6B6B6C6C6C4D4D2C4D6D8D6C6ACAAC8EC282400021210000;
defparam sp_inst_23.INIT_RAM_0E = 256'h37D58581D1B810690FF3D450CC8CAD8CADADADAD8C8CACACACACAC8C8C8C8CAC;
defparam sp_inst_23.INIT_RAM_0F = 256'h704C8EF12ED03555F0F011736F4C0F3052D0563A36104DEF6C8CC8A8ACCDCC6F;
defparam sp_inst_23.INIT_RAM_10 = 256'h969676765534559676B3D8F8CFAF14D3145619BB1CBEBEDB1AFA58D67491EECE;
defparam sp_inst_23.INIT_RAM_11 = 256'h05B43A97518F57FF7CFFFF5DBE3B993BBABA79375877732EE80D93D718B714B2;
defparam sp_inst_23.INIT_RAM_12 = 256'h618103A5A5E36140E2804750D2371131B0ADF0F26F0B2A8E2D103653128DAB2B;
defparam sp_inst_23.INIT_RAM_13 = 256'h8C8C6C6C6C6C4C4C4B6C8C2BC829CD52E3824000212101000021414141404040;
defparam sp_inst_23.INIT_RAM_14 = 256'hF4D4B2ED2B6CAD6BCCCCACACACADCDCCACACAC8C6B6B8BAC8C8CACACAC8C8C6C;
defparam sp_inst_23.INIT_RAM_15 = 256'h4FEED23C5D18D6337071B4902FF554908B8B8ACB0CCB6A8B4E725216B8536F6F;
defparam sp_inst_23.INIT_RAM_16 = 256'h769BB5EF13B59396FFFFDF7DBE1B79FBFADA3754D3D2F314B2D3D453F111108E;
defparam sp_inst_23.INIT_RAM_17 = 256'hBD3C5C7DFB7DBE1B7B5B1ADADABA59F7D60E67C8CF76D755763514557635F4D3;
defparam sp_inst_23.INIT_RAM_18 = 256'h2121A8AC70534E7252EFD4134B6E6F69AB892C0DB37330CDCA278C4E4E157D7E;
defparam sp_inst_23.INIT_RAM_19 = 256'h8BCCCD2B67A74B12E38220002141210000214140204040608181E26485E36140;
defparam sp_inst_23.INIT_RAM_1A = 256'h0CCCAB8CACADADAD8CACAC8C6B6B6B8B8CACCDEDEDCDAC8C4B4B4B4B4B4B4B4B;
defparam sp_inst_23.INIT_RAM_1B = 256'h4A6DAC08CFD9344AEC4EF06E2949AB49ECAFF0B08CAD5475D52F8B2A6CADADAC;
defparam sp_inst_23.INIT_RAM_1C = 256'hFDDDFEDDBCDDDD3BDA991795B61838D8F87BD91678F55192AE72F89F5EBBFB17;
defparam sp_inst_23.INIT_RAM_1D = 256'h5BFADA1B1BDADB3CDBDB376F094930189614149618B714B235D5AEF19BB68FD6;
defparam sp_inst_23.INIT_RAM_1E = 256'h32F398BAB956B0EFCBA96D0C8E6B8D73D38E2B8B15FE5D3E3B3BDA79DA3C5D7E;
defparam sp_inst_23.INIT_RAM_1F = 256'hE38220002141210121214120202040608160A16464E26140A0258611776F4E92;
defparam sp_inst_23.INIT_RAM_20 = 256'hCB8A8CEECD4B29496EAFCFAF6E0DCDAC4B4B2A0AEAEA0A0A8A8B8B4AA7A74C12;
defparam sp_inst_23.INIT_RAM_21 = 256'h77575634718D4C6CABAA89AB2FF417D7700E8C4A6A8ACACACCCCCCECCCACAC8C;
defparam sp_inst_23.INIT_RAM_22 = 256'hB6F73859799ABADBBABABA7A39F856B33193B8DC1D5D9E7DF98FCE749454B696;
defparam sp_inst_23.INIT_RAM_23 = 256'h7D1C1CBA1248C78DF4F83934D356B85775F27094B46F11F59DFEFFBE9E9E1C79;
defparam sp_inst_23.INIT_RAM_24 = 256'h5309EB90ACAB8F4E92D4F573B17196FC3C3C1BBA99DA3C5CDB1B5B5B5B5B7C9C;
defparam sp_inst_23.INIT_RAM_25 = 256'h01012141414140202080C143A5226060E284CC727151F2D236375817B5F55655;
defparam sp_inst_23.INIT_RAM_26 = 256'h3514F472B02EEDCDCDACAC8C8C8C8CACCB8B6B2AE8086CD1A161202020202100;
defparam sp_inst_23.INIT_RAM_27 = 256'hEE6B09ED349854AFAD8D6C6B8BCBEC0CECECECCCCCACAC8CEB8BACCD8C6A6EF3;
defparam sp_inst_23.INIT_RAM_28 = 256'hFB1CFBBB9A5AD85651F0F173B73D3CF77591F2116B6B74DAB43211D37675D250;
defparam sp_inst_23.INIT_RAM_29 = 256'h599634B639F8D5F29676107174D2957CDE9D7DBEDE5D9AF738599ABADBFB1C1C;
defparam sp_inst_23.INIT_RAM_2A = 256'h71B2D4D473B10FAE7518BA1B3C3CFBBA5C7D5CFAFA5B5BFA1BD9B52E8A4B8F51;
defparam sp_inst_23.INIT_RAM_2B = 256'hA2E30364A523606026C86A4928AE14147716549537738F31F6F1100F8C8F32EC;
defparam sp_inst_23.INIT_RAM_2C = 256'h6F909090909090908F0DAC8B6A8A2C0F8160200020202100210100000041A2C2;
defparam sp_inst_23.INIT_RAM_2D = 256'h2B4C8CACACCCEC0DCCCCCCACACACACACABCCAC8CEDF096DB5939B7D4F04E2E4E;
defparam sp_inst_23.INIT_RAM_2E = 256'hD3F0CC6BB0D8F73094F1D06E8A2D93B5906F6FD032B3359631302F2F104FECC8;
defparam sp_inst_23.INIT_RAM_2F = 256'hF7B310F354B71CFC9D5C7DBE7D7AF8F8BADBFB1C3C3C3C5D5C5D3D1CFCDB5AF8;
defparam sp_inst_23.INIT_RAM_30 = 256'h2C509558BAFB1C1C5C3B5C9D5CFB1B9DB8F44C474A5236D5D6759619D894308E;
defparam sp_inst_23.INIT_RAM_31 = 256'h86A7A7660831B7767437B95450F6F9720E73B876706F6F8B70919192B3D473D1;
defparam sp_inst_23.INIT_RAM_32 = 256'hB432D06F2DCCCC0C81612020200000000001416261402020204081E385640303;
defparam sp_inst_23.INIT_RAM_33 = 256'h8C8B8B8B8CACCCCD6BCCABCC729A5DDA9A7A183572F011527393B4B4D4D4D4B4;
defparam sp_inst_23.INIT_RAM_34 = 256'hF1D476D310F4F9DA38B12BEAED117373F65634CEA7430446C92B8CCDCDCCCDCD;
defparam sp_inst_23.INIT_RAM_35 = 256'h1B7DBE7D5996D79AFB1C3C5D3C3C3C5D5C7D5D3C3C1CBB593552EDC92AF0716D;
defparam sp_inst_23.INIT_RAM_36 = 256'h1A3B3B3C5C5C1BDA906BC9CC9377169455385977F2ADCB496B128F11B977373B;
defparam sp_inst_23.INIT_RAM_37 = 256'h74B591F35CFE5B9C78749090112FEDEDB012B0AD4C0F9292B5702B2B9158FBDB;
defparam sp_inst_23.INIT_RAM_38 = 256'hC2A161402000000000000020406181A1E324246507E785858141C3086E739433;
defparam sp_inst_23.INIT_RAM_39 = 256'h8C6BAC3159BE9DBADBDB79D735F435767697B7D8F8D8D8D8B77615B3116ECC8B;
defparam sp_inst_23.INIT_RAM_3A = 256'hBA99D6702B6CF277B977B20B25E1A2042687E94B6B8CACADAC8C8C8C8CACCCCD;
defparam sp_inst_23.INIT_RAM_3B = 256'h1C1C3C5D3C3C3C3C5C5D5D3C3C1CBB5A5631CDE9884A2C2CEE5356F4F43AFEDE;
defparam sp_inst_23.INIT_RAM_3C = 256'h4908CC5337F694B5BA3935904CAA28C7C6CA50333051D7B7BA3C3C39557639FC;
defparam sp_inst_23.INIT_RAM_3D = 256'hFF79710FB08EAE902EF1F1ED6BED502F7215F5D16C6CB1D61ABD7DFB5CFEB8AF;
defparam sp_inst_23.INIT_RAM_3E = 256'h2141414140202020218282C3658503E241C3A70DF1F29070532F759DFFFFFE1A;
defparam sp_inst_23.INIT_RAM_3F = 256'h5C1B9AF89696B7F839597A9A9A9A9A7A393918B7F4112EAC03E3A26120000000;

SP sp_inst_24 (
    .DO({sp_inst_24_dout_w[23:0],sp_inst_24_dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:8]})
);

defparam sp_inst_24.READ_MODE = 1'b0;
defparam sp_inst_24.WRITE_MODE = 2'b00;
defparam sp_inst_24.BIT_WIDTH = 8;
defparam sp_inst_24.BLK_SEL = 3'b001;
defparam sp_inst_24.RESET_MODE = "SYNC";
defparam sp_inst_24.INIT_RAM_00 = 256'h4A4A43434C4C443C080800000000000000000000000000000010213121000000;
defparam sp_inst_24.INIT_RAM_01 = 256'h424A525252524A4A5252524A4A4A4A4A4242424A4A4A4A4A4A4A4A4A524A4A4A;
defparam sp_inst_24.INIT_RAM_02 = 256'hBE5B7CAD9DC6D7B695859EA68D8D9E95CEDEEEFFFFC6753C242C3C5C6C5C4A3A;
defparam sp_inst_24.INIT_RAM_03 = 256'h3AB6BE746C7D95D7DEEFDEAD84524263DEE6E6F7EFB57B7CA5B68D748DB6CFAE;
defparam sp_inst_24.INIT_RAM_04 = 256'hC5B5A5A5A5ADBED7FFF6EEF6FFFFE6CEEEEEEEEEEEEEE6DEE6FEFED5BDE6C642;
defparam sp_inst_24.INIT_RAM_05 = 256'hBEADBE94638DAEB67522639DB695753B4BBEF6FEFEEFE7A5BEF7FFF7FFEFDEF7;
defparam sp_inst_24.INIT_RAM_06 = 256'h1008000000000000000000000000000000082129210800001821005BD6D6ADC6;
defparam sp_inst_24.INIT_RAM_07 = 256'h5252524A4A4A4A4A4A4A4A4A4A4A4A4A42424A4A4A4A4A4A52525A5353434343;
defparam sp_inst_24.INIT_RAM_08 = 256'h757D6D4C4454646DC5FFD5B3F6F79E5534446D756C4A42524A525A5A52524A4A;
defparam sp_inst_24.INIT_RAM_09 = 256'hE6F7E6C5AD73525B63628CB5835A739D9E6C64AEBE8C7C739DD7AD7CB6953B64;
defparam sp_inst_24.INIT_RAM_0A = 256'hD6E6EFE6DEE6F6FFEEEEF6EEEEE6EEF6DEDEE6FFEEA46B74B563529DC6C6D6EE;
defparam sp_inst_24.INIT_RAM_0B = 256'h5C43A6C695535C5C43E7FFF6FFC6ADBEFFE7FFFFEFF7F7C5FEFFFFDEA5847D85;
defparam sp_inst_24.INIT_RAM_0C = 256'h0000000000000000000819292108000008090095D6CEB5A58DAEA58DB6CF967D;
defparam sp_inst_24.INIT_RAM_0D = 256'h52524A4A4A4A4A4A42424A4A4A4A4A4A5A5A5A524A425B6C1810000000000000;
defparam sp_inst_24.INIT_RAM_0E = 256'hEFEE7259DDF79E4C658595744A4A525252525A5A5A525252525252524A4A4A52;
defparam sp_inst_24.INIT_RAM_0F = 256'h8C6B73836B739D9D646C7D957C6384848D7CB6D7AE7D5C6C4C442B23444C4C65;
defparam sp_inst_24.INIT_RAM_10 = 256'hEEEEEEE6E6DEE6EED6C5E6E69C8CAE9D9DB5D6E6E7F7FFF6EFEED6C5B5947B7B;
defparam sp_inst_24.INIT_RAM_11 = 256'h1AA5EFDEAD84BEFFE7FFFFF7FFEFD6EFE6E6DED6D6D6B58C4A74ADDEF7F6EEE5;
defparam sp_inst_24.INIT_RAM_12 = 256'h000011212110000808002A6C94C695958D6C8484745C5475755CA6A68D746C43;
defparam sp_inst_24.INIT_RAM_13 = 256'h4A4A4A4242424242424A524A393A639518100000000000000000000000000000;
defparam sp_inst_24.INIT_RAM_14 = 256'h9D9D8452424A52425A5A5A5A5A5A5A5252525252525252524A52525252524A4A;
defparam sp_inst_24.INIT_RAM_15 = 256'h746B94EFF7C6BDA58D8DA58474A59E7D4C4C44444D443C448DBEC6E7F7B68575;
defparam sp_inst_24.INIT_RAM_16 = 256'hDEFFBD7395ADA5C6F7FFFFFFF7E7D6F6EEE6CEB5A4A4A4AD9CA4A49483847C63;
defparam sp_inst_24.INIT_RAM_17 = 256'hEFE7F7F7EEF7FFE7E7E7DFE6EEEEEEE5BD7C42529CD6EEE6EEDEDEE6E6DED5D5;
defparam sp_inst_24.INIT_RAM_18 = 256'h09012A5384A57C95A684AD95536C7D546C2A546D8DA6A6633A326B7C74AEEFFF;
defparam sp_inst_24.INIT_RAM_19 = 256'h3A424A4229295B8D181000000000000000000000000000000000001919100808;
defparam sp_inst_24.INIT_RAM_1A = 256'h5B5A5A5A5A5A525252525A525252525A4A52525A5A52524A424242423A3A3A3A;
defparam sp_inst_24.INIT_RAM_1B = 256'h64746B3A73C6A654646D755D3434443C64859595746C9696A5744A4252524A4A;
defparam sp_inst_24.INIT_RAM_1C = 256'hE7EFFFFFEFEFF7EFE6DEC6BDC5CED6CDCDE6CDBDBDAC8C8C83A4D5FFFFDEDEB6;
defparam sp_inst_24.INIT_RAM_1D = 256'hEFE6DEEFEFDEDEEFEEE6C68C535BA5E7EEDEDEEEFFF6DECDE6CD7373C6AD8CDE;
defparam sp_inst_24.INIT_RAM_1E = 256'hAEADCED6CEB68D8D742A5C655C5C8D9D845B535BA6F7F7FFE7E7DEDEE6EFEFEF;
defparam sp_inst_24.INIT_RAM_1F = 256'h181000000008000000000000000000000000001119100808001A227DBE847C95;
defparam sp_inst_24.INIT_RAM_20 = 256'h5A525A6262524A52737B7B7B736B625A4A4A4A42414142424A4A4A4229295B95;
defparam sp_inst_24.INIT_RAM_21 = 256'hC6BEB6A6855C4C4C2C2C34548DB5AE9D635B4A424A525A5A6262625A5A5A524A;
defparam sp_inst_24.INIT_RAM_22 = 256'hBDC5CED6D6DEDEE6DEE6DEDED6C5B5A4949CC5E6EFF7FFF7DD8B7BA5A59DB5B5;
defparam sp_inst_24.INIT_RAM_23 = 256'hEFE7EFE6A55B537DD5FEFFEEDDEEF6DEB59C8CADAD8C9DC5F7FFFFFFF7F7E7D6;
defparam sp_inst_24.INIT_RAM_24 = 256'hA54B4B6D545C8D959DADB5A5948CB5DEEFF7EFDEDEE6F7F7E6EFF7F7EFEFF7FF;
defparam sp_inst_24.INIT_RAM_25 = 256'h0000000000000000000000112119081010195B8D8D95A5ADC6C6C6C6B5BDC6C6;
defparam sp_inst_24.INIT_RAM_26 = 256'hADADA4947B6B62625A5A5A5A5A5A5A5A5A524A42313A638C1008000000000000;
defparam sp_inst_24.INIT_RAM_27 = 256'h5C443C64AECEA5634A4A42424A525A636262625A5A52524A5A525A625A527BA4;
defparam sp_inst_24.INIT_RAM_28 = 256'hEEEFEEE6DED6C5B594838394BDEFEFC5BD94948553539DCEAD9D8D9DAEA68D75;
defparam sp_inst_24.INIT_RAM_29 = 256'hFFEEE6F6FFEEC5A4B5B5848CAD9CBDFFFFF7F7FFFFEFD6C5CED6D6DEE6E6E7EF;
defparam sp_inst_24.INIT_RAM_2A = 256'h959DA5AD9D8C7C73B5CEDEEFF7F7EEE6F7F7EFE6E6EFEFE6F7DEAD745B74A5C6;
defparam sp_inst_24.INIT_RAM_2B = 256'h08080911211108082A3A4B43437CB6B6CEBEADB5C6AD94A5B58C7D755C7D9E74;
defparam sp_inst_24.INIT_RAM_2C = 256'h7B7B7B7B7B7B7B7B7B6B5A524A4A637C10080000000000000000000000000808;
defparam sp_inst_24.INIT_RAM_2D = 256'h42424A52525A5A635A5A5A5A525252525A5A5A5A628BBDE6D6CEBDA483736B73;
defparam sp_inst_24.INIT_RAM_2E = 256'hA48362527BC5C58CA58C7C6C4B6C9DAD84848484959DA6B695856D75857C5A31;
defparam sp_inst_24.INIT_RAM_2F = 256'hBD947C9CADC5F7F6F7EFF7FFF7D6C5C5DEDEE6EFEFEFEFEFF7F7F7EFEEE6D6C5;
defparam sp_inst_24.INIT_RAM_30 = 256'h6B8CB5D6E6EEF7F7EFEFF7F7F7E6EFF7EEBD6C3B64BEFFFEF6E6EEF7E6B57C5B;
defparam sp_inst_24.INIT_RAM_31 = 256'h3232322A4395C6C6ADC6D6AD8CBDDEAD7CA5CEB68D7D7554858D95959DA59D8C;
defparam sp_inst_24.INIT_RAM_32 = 256'hA49483736B5A5A63100800000000000000000008000000000000000821211119;
defparam sp_inst_24.INIT_RAM_33 = 256'h525252525252525A525A5A6294DEF7E6DED6C6AD94838C949C9CA4A4A4A4A4A4;
defparam sp_inst_24.INIT_RAM_34 = 256'h8CA5B69D8DADD6DEC6945B527395A5A5C5B68E5C2A11192131424A525252525A;
defparam sp_inst_24.INIT_RAM_35 = 256'hE7F7FFF7CEB5BDD6E6E7EFEFEFEFEFEFEFF7EFEFEFEFDECEAD8C62414A839473;
defparam sp_inst_24.INIT_RAM_36 = 256'hE7EFEFEFEFEFE7DEAD7C6384C6F7FFFEE6FFFFD6945B3A22538D748DCECECEEF;
defparam sp_inst_24.INIT_RAM_37 = 256'hADB594A4EFFFE7EFCEB59C949585645C85968564647D9D9DB58C636394D6EEE6;
defparam sp_inst_24.INIT_RAM_38 = 256'h10100800000000000000000000000808101919213231212101011143749DADA5;
defparam sp_inst_24.INIT_RAM_39 = 256'h52525A8CD6FFFFDEE6DED6BDADA4ADB5BDBDC5C5CDCDC5C5C5BDADA48C735A52;
defparam sp_inst_24.INIT_RAM_3A = 256'hD6D6BD8C636B9CCEDEB67D3C0A000011212939424A4A4A525252525252525A5A;
defparam sp_inst_24.INIT_RAM_3B = 256'hE7EFEFEFEFEFEFEFEFF7EFEFEFEFDED6AD845A41314A6B6373A5BEB5BDE7FFFF;
defparam sp_inst_24.INIT_RAM_3C = 256'h5C649CE6FFFEEEEEFFFFCE8C533222112A4B7D9E8595CECEDEEFEFCEADB5CEE6;
defparam sp_inst_24.INIT_RAM_3D = 256'hFFDE9C94947C6C757D8D8564546C85859DAEB58C6B6B9CC5DFF7F7DEEFFFD694;
defparam sp_inst_24.INIT_RAM_3E = 256'h0000000000000000000808102929191001113A6C949C8C8CAD8CB5F7FFFFFFE7;
defparam sp_inst_24.INIT_RAM_3F = 256'hEFE7D6C5BDB5BDC5CED6D6DEDEDEDED6D6CECEBDA4846B5A1918100800000000;

SP sp_inst_25 (
    .DO({sp_inst_25_dout_w[15:0],sp_inst_25_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_9}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_25.READ_MODE = 1'b0;
defparam sp_inst_25.WRITE_MODE = 2'b00;
defparam sp_inst_25.BIT_WIDTH = 16;
defparam sp_inst_25.BLK_SEL = 3'b001;
defparam sp_inst_25.RESET_MODE = "SYNC";
defparam sp_inst_25.INIT_RAM_00 = 256'h4AAD4AAD4A8C528C52AC52AC52AC5AAC62EE4A2A6B2DC5D7F77DEF3BE6FBF77D;
defparam sp_inst_25.INIT_RAM_01 = 256'hBE169DD46D51440C1A66010200610081086210A31904296631A83A09424B4A6C;
defparam sp_inst_25.INIT_RAM_02 = 256'h62EB9470B594C5F6DEB9FF9DFF9DF6FBFFDFFFBEE6FBC618B575AD75BDD6BDF6;
defparam sp_inst_25.INIT_RAM_03 = 256'hEF5CEF5CEF5DEF3CEF3CE71CDEBBCE39B5B77BD04A6B39C9318739C84A6A5ACA;
defparam sp_inst_25.INIT_RAM_04 = 256'hCE58CE38B5769C929CB3BDB7D67ADEBBE6FBEF1CEF3CEF3CEF3CEF3CEF3CEF3C;
defparam sp_inst_25.INIT_RAM_05 = 256'hF719BD937BED52EA3A6932483AAA536D6CAD95F274CD6CAD95B18D509D51BE35;
defparam sp_inst_25.INIT_RAM_06 = 256'h94B0A553D6BAFFDEE75BAD737C2C73EA6C8AA5AFEED5FEF6FE96FE96F718EFB9;
defparam sp_inst_25.INIT_RAM_07 = 256'h74CD856F7D906D4E6D6E85F18DF17D6F855095B1A5F3AE34ADF49D73844F634B;
defparam sp_inst_25.INIT_RAM_08 = 256'hA512F77CFFFFFFDFFFFFFFBEEF3CFFDED699EF3CF73BDE79C5F6A5738D118D51;
defparam sp_inst_25.INIT_RAM_09 = 256'h31A641E739C641C64A4842272964190219A44B096BCC6BAC7BED842F94B1AD53;
defparam sp_inst_25.INIT_RAM_0A = 256'h2124210318E310820041000000000000002000200000000008201040108118A2;
defparam sp_inst_25.INIT_RAM_0B = 256'hDEBADEBADEDBDEDBDEDBDEDBDEDBDEDADE9BD67AD679C618B59694B373B05AEE;
defparam sp_inst_25.INIT_RAM_0C = 256'h5AAD5AAC8C31D699F79DE6DAE6DAFFBDF75CE6FBD659C5D7BDB6BDD7CE19CE59;
defparam sp_inst_25.INIT_RAM_0D = 256'h088108610861088210E4214629A829C83A2B3A2B424B426B4A8C528C528C52AC;
defparam sp_inst_25.INIT_RAM_0E = 256'hE6DCFF9FFFDFE6FBB595A513B595C6589D738D7275515C4E42A82123108110A1;
defparam sp_inst_25.INIT_RAM_0F = 256'hA5156B2E39E93188318741E95AEC738E738EBDB6F75CF77CEEFADEBAE6BAEF1C;
defparam sp_inst_25.INIT_RAM_10 = 256'hDEBAE6DBE71CE71CE71CE71CE71CEF1CE73CEF3CE73CE71CE6FCDEDBCE59BDD7;
defparam sp_inst_25.INIT_RAM_11 = 256'hCEB7B5F495119D72A593A573AD749470AD3494927BAF738E8C31AD56CE19D67A;
defparam sp_inst_25.INIT_RAM_12 = 256'hD612F716FF78FF17FED7FF18F739E6F9AD12947073CE636D5B6C6BCD84B09D52;
defparam sp_inst_25.INIT_RAM_13 = 256'h750D7D4E856F8D708D719D929D929D72634B632B9491CE58A55252E75B059D2C;
defparam sp_inst_25.INIT_RAM_14 = 256'hEF3CEF3BE6DADEB9EF3BEF5BC617947084AE850F752F64ED5CED654E650E64AC;
defparam sp_inst_25.INIT_RAM_15 = 256'h320752CA5ACA62CA734C7BCD9CD0C656FFFEEF3BF77DFFFFFFFFEF5DF77DF77D;
defparam sp_inst_25.INIT_RAM_16 = 256'h00000000000018823986730C9C91BD75D678DE99D617C595BD749CB16B6B52A8;
defparam sp_inst_25.INIT_RAM_17 = 256'hE6DCD6BBCE79C637B5D79D147BF15AEE2103190318C310820041000000210021;
defparam sp_inst_25.INIT_RAM_18 = 256'hF77DE6DACE38BDB6BDD7CE39D69ADEDBDEFBDEFBDEFBDEFBDEFBDEFBDEDBDEDB;
defparam sp_inst_25.INIT_RAM_19 = 256'h2168298931C93A0A424B4A6B528B528C4A4B6B4FA4F4D679EF5BF77CEF3BEF1B;
defparam sp_inst_25.INIT_RAM_1A = 256'h9D93853174AF6C0E630B520741853964212318C108600020006108A310E410E5;
defparam sp_inst_25.INIT_RAM_1B = 256'hCE59DEBAD699CE58D699CE79BDD7B5B6E6BBE6DCD65AB5769CB294B294F29D13;
defparam sp_inst_25.INIT_RAM_1C = 256'hDEFBE71BE71BDEFBDEDBD69AC618B57673B0528B31A82967318852AC8C51AD55;
defparam sp_inst_25.INIT_RAM_1D = 256'h84106B4D62CB6B2D83D09493B597D67BD679DE9ADEDBE6DBE6DBE6DBE6FBE6FB;
defparam sp_inst_25.INIT_RAM_1E = 256'h9CD2AD55A55594F3A595CEB9D6B7B5B3A4B2C5D6C5D6CE58CE59AD14A493A493;
defparam sp_inst_25.INIT_RAM_1F = 256'hBE16A553842F6B6C636A846CB60FDF53FF19FED7F6B5EF16F7B9F77AD616B4B2;
defparam sp_inst_25.INIT_RAM_20 = 256'h73CC7CAE7D2F6D4F5D0D5D0D650D650D64EB6D2C754E7D4E8570957195719551;
defparam sp_inst_25.INIT_RAM_21 = 256'hD677FFBDFFDEE6FCEF1CFF9EF75DE6DBF75CE6FBE71BEF5CEF7CEEFBCDB69BEF;
defparam sp_inst_25.INIT_RAM_22 = 256'hDE79EEDAEE99E658E678CDF69CD07C0D738E5ACB5269838EACF29CB0A532E739;
defparam sp_inst_25.INIT_RAM_23 = 256'h18E318E310C208820041002000210841000028E462EBA4D3D638EEDAEEDBEEBA;
defparam sp_inst_25.INIT_RAM_24 = 256'hDEDBE6FBE6FBE6FBE6FBE6FBE6FBDEDBDEFBDEFBDEDBCE59BDD7A4F47BD05AEC;
defparam sp_inst_25.INIT_RAM_25 = 256'h4A8C632E9CD3CE38DE99E6DAEF3BE73BEF3DC618B597BDD7C5F8CE39DEBBDEBB;
defparam sp_inst_25.INIT_RAM_26 = 256'h41E8210408410840088108810060008010E310E31924298731C839E9422B4A8C;
defparam sp_inst_25.INIT_RAM_27 = 256'hC5F7C5F7BDD7B596B575BDB6BDB6BDB69D348C9294919CF29CD18C2F736C5A69;
defparam sp_inst_25.INIT_RAM_28 = 256'h4A8C31C9212618A349E883CEACF2DE98EF3BE71BE6FBE6FBDEDAD699CE18BDD7;
defparam sp_inst_25.INIT_RAM_29 = 256'hBD96C5D7D639DE7ADE9ADE9ADE9ADE9ADE9BDEBBDE9BD65AC619B577949373B0;
defparam sp_inst_25.INIT_RAM_2A = 256'hAD94B5B6C639B6578D92750E84CF846F6BAE52EB42494A6B52AC630E8411A515;
defparam sp_inst_25.INIT_RAM_2B = 256'hF6F7E675FF18FF7ADE57BD94BDB5B595EF7EC678ADF4B634B634BE55BDF6AD75;
defparam sp_inst_25.INIT_RAM_2C = 256'h74CF855095D17D2E7D6D54894CCA550B750D858E95AFA591AD73CDB4EE76FF16;
defparam sp_inst_25.INIT_RAM_2D = 256'hEF7CEF3CF77DEF1CB595846E748C7D2D85D16D2E5CCB54AB64CC856F8D507C4D;
defparam sp_inst_25.INIT_RAM_2E = 256'h6B4D632C632C5ACB6B2B8C0EACD0E676AD14E6DAE6FBDEDAE6DAE6FBEF7DEF5C;
defparam sp_inst_25.INIT_RAM_2F = 256'h838EACF3D658E6DAE6DADEDADEDADEDAE6DADEBAE6DBE6BAD659CE18B53483CF;
defparam sp_inst_25.INIT_RAM_30 = 256'hDEDBDEDBD6BACE59B5B79CF47BAF5ACC108110A208A200210041000000002903;
defparam sp_inst_25.INIT_RAM_31 = 256'hD69BB596AD35B597BDD8CE39DEBBDEBBDEDBE6FBE6FBE6FBE6FBE6FBE6FBDEDB;
defparam sp_inst_25.INIT_RAM_32 = 256'h0061006208A319052146298831C9422B422B5ACD8C72C5D7CE38D678DEDADEDA;
defparam sp_inst_25.INIT_RAM_33 = 256'hAD9694D394D2AD74B5B5B5549450732C41E82104084108400881088100600080;
defparam sp_inst_25.INIT_RAM_34 = 256'hF77CEF5CEF3BE71BE6FBDEBAD659C618C618CE38C617BDD7BDB6C5F7C5F7BDD7;
defparam sp_inst_25.INIT_RAM_35 = 256'hBD97BD97B576AD159CB483F15AED4209298821262126312562ABA492C595EEFA;
defparam sp_inst_25.INIT_RAM_36 = 256'h5B2C426931C839E93A0A422A5AED7BD08BF09431A4B3AD14B555BD76BD96BD96;
defparam sp_inst_25.INIT_RAM_37 = 256'hA5357C0F6BEC84CE9D50A592AD95AD55BDF6BDD7BE18A5B56CAE4C0A53CA5B4B;
defparam sp_inst_25.INIT_RAM_38 = 256'h64EB6D0C7D0C8D0FA531C594DE14EE94FF17EEB6F718EEF8C5B4BD94D678DEB9;
defparam sp_inst_25.INIT_RAM_39 = 256'h7D6F6D2E650C5CEC64EC85909DB2951085318D929E12856E858E5CAA54CA550B;
defparam sp_inst_25.INIT_RAM_3A = 256'h9C91D658DEBADEBADEDAE6FBF77DEF5CF79DEF3CDE7AA4D36B6C63AB7CEE8DAF;
defparam sp_inst_25.INIT_RAM_3B = 256'hE6FBE6DAE6FBE6DADE79CE38B5548BEF632C5ACB528A31A639A54A06628793EC;
defparam sp_inst_25.INIT_RAM_3C = 256'h0860004000610000004108622104736DC5B6D658E6BADEBADE99DEBAE6DADEFA;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce_w)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(spx9_inst_0_dout[0]),
  .I1(spx9_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(spx9_inst_2_dout[0]),
  .I1(spx9_inst_3_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(spx9_inst_4_dout[0]),
  .I1(spx9_inst_5_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(spx9_inst_6_dout[0]),
  .I1(spx9_inst_7_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(sp_inst_23_dout[0]),
  .I1(sp_inst_25_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(mux_o_11),
  .I1(mux_o_12),
  .S0(dff_q_2)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_13),
  .I1(mux_o_14),
  .S0(dff_q_2)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(mux_o_17),
  .I1(mux_o_18),
  .S0(dff_q_1)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(sp_inst_15_dout[0]),
  .I1(mux_o_16),
  .S0(dff_q_1)
);
MUX2 mux_inst_23 (
  .O(dout[0]),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(spx9_inst_0_dout[1]),
  .I1(spx9_inst_1_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(spx9_inst_2_dout[1]),
  .I1(spx9_inst_3_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(spx9_inst_4_dout[1]),
  .I1(spx9_inst_5_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(spx9_inst_6_dout[1]),
  .I1(spx9_inst_7_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(sp_inst_23_dout[1]),
  .I1(sp_inst_25_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_2)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_37),
  .I1(mux_o_38),
  .S0(dff_q_2)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(mux_o_41),
  .I1(mux_o_42),
  .S0(dff_q_1)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sp_inst_15_dout[1]),
  .I1(mux_o_40),
  .S0(dff_q_1)
);
MUX2 mux_inst_47 (
  .O(dout[1]),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_0)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(spx9_inst_0_dout[2]),
  .I1(spx9_inst_1_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(spx9_inst_2_dout[2]),
  .I1(spx9_inst_3_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(spx9_inst_4_dout[2]),
  .I1(spx9_inst_5_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(spx9_inst_6_dout[2]),
  .I1(spx9_inst_7_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(sp_inst_23_dout[2]),
  .I1(sp_inst_25_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(mux_o_59),
  .I1(mux_o_60),
  .S0(dff_q_2)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(mux_o_61),
  .I1(mux_o_62),
  .S0(dff_q_2)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_65),
  .I1(mux_o_66),
  .S0(dff_q_1)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(sp_inst_16_dout[2]),
  .I1(mux_o_64),
  .S0(dff_q_1)
);
MUX2 mux_inst_71 (
  .O(dout[2]),
  .I0(mux_o_69),
  .I1(mux_o_70),
  .S0(dff_q_0)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(spx9_inst_0_dout[3]),
  .I1(spx9_inst_1_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(spx9_inst_2_dout[3]),
  .I1(spx9_inst_3_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(spx9_inst_4_dout[3]),
  .I1(spx9_inst_5_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(spx9_inst_6_dout[3]),
  .I1(spx9_inst_7_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(sp_inst_23_dout[3]),
  .I1(sp_inst_25_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_2)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_2)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_89),
  .I1(mux_o_90),
  .S0(dff_q_1)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(sp_inst_16_dout[3]),
  .I1(mux_o_88),
  .S0(dff_q_1)
);
MUX2 mux_inst_95 (
  .O(dout[3]),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(dff_q_0)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(spx9_inst_0_dout[4]),
  .I1(spx9_inst_1_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(spx9_inst_2_dout[4]),
  .I1(spx9_inst_3_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(spx9_inst_4_dout[4]),
  .I1(spx9_inst_5_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(spx9_inst_6_dout[4]),
  .I1(spx9_inst_7_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(sp_inst_23_dout[4]),
  .I1(sp_inst_25_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_2)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_2)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(dff_q_1)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(sp_inst_17_dout[4]),
  .I1(mux_o_112),
  .S0(dff_q_1)
);
MUX2 mux_inst_119 (
  .O(dout[4]),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_0)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(spx9_inst_0_dout[5]),
  .I1(spx9_inst_1_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(spx9_inst_2_dout[5]),
  .I1(spx9_inst_3_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(spx9_inst_4_dout[5]),
  .I1(spx9_inst_5_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(spx9_inst_6_dout[5]),
  .I1(spx9_inst_7_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sp_inst_23_dout[5]),
  .I1(sp_inst_25_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(mux_o_131),
  .I1(mux_o_132),
  .S0(dff_q_2)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(dff_q_2)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_1)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(sp_inst_17_dout[5]),
  .I1(mux_o_136),
  .S0(dff_q_1)
);
MUX2 mux_inst_143 (
  .O(dout[5]),
  .I0(mux_o_141),
  .I1(mux_o_142),
  .S0(dff_q_0)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(spx9_inst_0_dout[6]),
  .I1(spx9_inst_1_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(spx9_inst_2_dout[6]),
  .I1(spx9_inst_3_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(spx9_inst_4_dout[6]),
  .I1(spx9_inst_5_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(spx9_inst_6_dout[6]),
  .I1(spx9_inst_7_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(sp_inst_23_dout[6]),
  .I1(sp_inst_25_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_155),
  .I1(mux_o_156),
  .S0(dff_q_2)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_157),
  .I1(mux_o_158),
  .S0(dff_q_2)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(dff_q_1)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(sp_inst_18_dout[6]),
  .I1(mux_o_160),
  .S0(dff_q_1)
);
MUX2 mux_inst_167 (
  .O(dout[6]),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_0)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(spx9_inst_0_dout[7]),
  .I1(spx9_inst_1_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(spx9_inst_2_dout[7]),
  .I1(spx9_inst_3_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(spx9_inst_4_dout[7]),
  .I1(spx9_inst_5_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(spx9_inst_6_dout[7]),
  .I1(spx9_inst_7_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(sp_inst_23_dout[7]),
  .I1(sp_inst_25_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_2)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_2)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(mux_o_185),
  .I1(mux_o_186),
  .S0(dff_q_1)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(sp_inst_18_dout[7]),
  .I1(mux_o_184),
  .S0(dff_q_1)
);
MUX2 mux_inst_191 (
  .O(dout[7]),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_0)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(spx9_inst_0_dout[8]),
  .I1(spx9_inst_1_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(spx9_inst_2_dout[8]),
  .I1(spx9_inst_3_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(spx9_inst_4_dout[8]),
  .I1(spx9_inst_5_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(spx9_inst_6_dout[8]),
  .I1(spx9_inst_7_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(sp_inst_24_dout[8]),
  .I1(sp_inst_25_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_2)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_2)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(mux_o_209),
  .I1(mux_o_210),
  .S0(dff_q_1)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(sp_inst_19_dout[8]),
  .I1(mux_o_208),
  .S0(dff_q_1)
);
MUX2 mux_inst_215 (
  .O(dout[8]),
  .I0(mux_o_213),
  .I1(mux_o_214),
  .S0(dff_q_0)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(sp_inst_24_dout[9]),
  .I1(sp_inst_25_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(sp_inst_19_dout[9]),
  .I1(mux_o_222),
  .S0(dff_q_1)
);
MUX2 mux_inst_228 (
  .O(dout[9]),
  .I0(sp_inst_8_dout[9]),
  .I1(mux_o_227),
  .S0(dff_q_0)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(sp_inst_24_dout[10]),
  .I1(sp_inst_25_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(sp_inst_20_dout[10]),
  .I1(mux_o_235),
  .S0(dff_q_1)
);
MUX2 mux_inst_241 (
  .O(dout[10]),
  .I0(sp_inst_9_dout[10]),
  .I1(mux_o_240),
  .S0(dff_q_0)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(sp_inst_24_dout[11]),
  .I1(sp_inst_25_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(sp_inst_20_dout[11]),
  .I1(mux_o_248),
  .S0(dff_q_1)
);
MUX2 mux_inst_254 (
  .O(dout[11]),
  .I0(sp_inst_10_dout[11]),
  .I1(mux_o_253),
  .S0(dff_q_0)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(sp_inst_24_dout[12]),
  .I1(sp_inst_25_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(sp_inst_21_dout[12]),
  .I1(mux_o_261),
  .S0(dff_q_1)
);
MUX2 mux_inst_267 (
  .O(dout[12]),
  .I0(sp_inst_11_dout[12]),
  .I1(mux_o_266),
  .S0(dff_q_0)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(sp_inst_24_dout[13]),
  .I1(sp_inst_25_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(sp_inst_21_dout[13]),
  .I1(mux_o_274),
  .S0(dff_q_1)
);
MUX2 mux_inst_280 (
  .O(dout[13]),
  .I0(sp_inst_12_dout[13]),
  .I1(mux_o_279),
  .S0(dff_q_0)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(sp_inst_24_dout[14]),
  .I1(sp_inst_25_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(sp_inst_22_dout[14]),
  .I1(mux_o_287),
  .S0(dff_q_1)
);
MUX2 mux_inst_293 (
  .O(dout[14]),
  .I0(sp_inst_13_dout[14]),
  .I1(mux_o_292),
  .S0(dff_q_0)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(sp_inst_24_dout[15]),
  .I1(sp_inst_25_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(sp_inst_22_dout[15]),
  .I1(mux_o_300),
  .S0(dff_q_1)
);
MUX2 mux_inst_306 (
  .O(dout[15]),
  .I0(sp_inst_14_dout[15]),
  .I1(mux_o_305),
  .S0(dff_q_0)
);
endmodule //Gowin_SP
